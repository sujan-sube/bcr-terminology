C0006142|T047|dctl adenoca|breast cancer_C0006142
C0006142|T047|lobular adenocarcinoma|breast cancer_C0006142
C0006142|T047|breast carcinoma|breast cancer_C0006142
C0006142|T047|ca br|breast cancer_C0006142
C0006142|T047|adenocarc lobular|breast cancer_C0006142
C0006142|T047|ca breast|breast cancer_C0006142
C0006142|T047|ca dctl|breast cancer_C0006142
C0006142|T047|breast carc|breast cancer_C0006142
C0006142|T047|ca ductal|breast cancer_C0006142
C0006142|T047|adenocarc ductal|breast cancer_C0006142
C0006142|T047|adenocarc dctl|breast cancer_C0006142
C0006142|T047|adenocarc breast|breast cancer_C0006142
C0006142|T047|adenocarc br|breast cancer_C0006142
C0006142|T047|cancer br|breast cancer_C0006142
C0006142|T047|lobular ca|breast cancer_C0006142
C0006142|T047|ca lobular|breast cancer_C0006142
C0006142|T047|breast cancer|breast cancer_C0006142
C0006142|T047|breast ca|breast cancer_C0006142
C0006142|T047|breast adenocarcinoma|breast cancer_C0006142
C0006142|T047|adenocarcinoma breast|breast cancer_C0006142
C0006142|T047|adenocarcinoma dctl|breast cancer_C0006142
C0006142|T047|adenocarcinoma ductal|breast cancer_C0006142
C0006142|T047|adenocarcinoma lobular|breast cancer_C0006142
C0006142|T047|br adenoca|breast cancer_C0006142
C0006142|T047|br adenocarc|breast cancer_C0006142
C0006142|T047|br adenocarcinoma|breast cancer_C0006142
C0006142|T047|br ca|breast cancer_C0006142
C0006142|T047|br cancer|breast cancer_C0006142
C0006142|T047|lobular adenoca|breast cancer_C0006142
C0006142|T047|br carc|breast cancer_C0006142
C0006142|T047|br carcinoma|breast cancer_C0006142
C0006142|T047|breast adenoca|breast cancer_C0006142
C0006142|T047|breast adenocarc|breast cancer_C0006142
C0006142|T047|lobular adenocarc|breast cancer_C0006142
C0006142|T047|adenocarcinoma br|breast cancer_C0006142
C0006142|T047|cancer dctl|breast cancer_C0006142
C0006142|T047|cancer breast|breast cancer_C0006142
C0006142|T047|cancer lobular|breast cancer_C0006142
C0006142|T047|carcinoma br|breast cancer_C0006142
C0006142|T047|carcinoma breast|breast cancer_C0006142
C0006142|T047|carcinoma dctl|breast cancer_C0006142
C0006142|T047|carcinoma ductal|breast cancer_C0006142
C0006142|T047|carcinoma lobular|breast cancer_C0006142
C0006142|T047|dctl carc|breast cancer_C0006142
C0006142|T047|adenoca lobular|breast cancer_C0006142
C0006142|T047|dctl cancer|breast cancer_C0006142
C0006142|T047|dctl ca|breast cancer_C0006142
C0006142|T047|dctl adenocarcinoma|breast cancer_C0006142
C0006142|T047|dctl adenocarc|breast cancer_C0006142
C0006142|T047|adenoca ductal|breast cancer_C0006142
C0006142|T047|adenoca dctl|breast cancer_C0006142
C0006142|T047|adenoca breast|breast cancer_C0006142
C0006142|T047|adenoca br|breast cancer_C0006142
C0006142|T047|dctl carcinoma|breast cancer_C0006142
C0006142|T047|cancer ductal|breast cancer_C0006142
C0006142|T047|ductal adenoca|breast cancer_C0006142
C0006142|T047|ductal adenocarcinoma|breast cancer_C0006142
C0006142|T047|lobular cancer|breast cancer_C0006142
C0006142|T047|ductal carcinoma|breast cancer_C0006142
C0006142|T047|ductal carc|breast cancer_C0006142
C0006142|T047|carc br|breast cancer_C0006142
C0006142|T047|lobular carc|breast cancer_C0006142
C0006142|T047|ductal adenocarc|breast cancer_C0006142
C0006142|T047|carc dctl|breast cancer_C0006142
C0006142|T047|carc breast|breast cancer_C0006142
C0006142|T047|carc lobular|breast cancer_C0006142
C0006142|T047|lobular carcinoma|breast cancer_C0006142
C0006142|T047|ductal cancer|breast cancer_C0006142
C0006142|T047|ductal ca|breast cancer_C0006142
C0006142|T047|carc ductal|breast cancer_C0006142
C0007097|T047|carc|cancer_C0007097
C0007097|T047|ca|cancer_C0007097
C0007097|T047|cancer|cancer_C0007097
C0007097|T047|carcinoma|cancer_C0007097
C0007097|T047|adenocarcinoma|cancer_C0007097
C0007097|T047|adenoca|cancer_C0007097
C0007097|T047|adenocarc|cancer_C0007097
C0007099|T047|in-situ carcinoma|intraductal cancer_C0007099
C0007099|T047|intraductl adenocarc|intraductal cancer_C0007099
C0007099|T047|carc intraductl|intraductal cancer_C0007099
C0007099|T047|in situ adenoca|intraductal cancer_C0007099
C0007099|T047|carcinoma intraductl|intraductal cancer_C0007099
C0007099|T047|carcinoma intraductal|intraductal cancer_C0007099
C0007099|T047|intraductl adenoca|intraductal cancer_C0007099
C0007099|T047|carcinoma in-situ|intraductal cancer_C0007099
C0007099|T047|carcinoma in situ|intraductal cancer_C0007099
C0007099|T047|intraductal cancer|intraductal cancer_C0007099
C0007099|T047|intraductal adenocarc|intraductal cancer_C0007099
C0007099|T047|intraductal adenoca|intraductal cancer_C0007099
C0007099|T047|in-situ adenoca|intraductal cancer_C0007099
C0007099|T047|in situ ca|intraductal cancer_C0007099
C0007099|T047|intraductal carc|intraductal cancer_C0007099
C0007099|T047|intraductal adenocarcinoma|intraductal cancer_C0007099
C0007099|T047|in situ carcinoma|intraductal cancer_C0007099
C0007099|T047|cancer intraductl|intraductal cancer_C0007099
C0007099|T047|cancer intraductal|intraductal cancer_C0007099
C0007099|T047|cancer in-situ|intraductal cancer_C0007099
C0007099|T047|intraductal carcinoma|intraductal cancer_C0007099
C0007099|T047|in situ carc|intraductal cancer_C0007099
C0007099|T047|cancer in situ|intraductal cancer_C0007099
C0007099|T047|in situ cancer|intraductal cancer_C0007099
C0007099|T047|carc in situ|intraductal cancer_C0007099
C0007099|T047|carc in-situ|intraductal cancer_C0007099
C0007099|T047|carc intraductal|intraductal cancer_C0007099
C0007099|T047|adenocarc in situ|intraductal cancer_C0007099
C0007099|T047|ca intraductl|intraductal cancer_C0007099
C0007099|T047|in-situ adenocarc|intraductal cancer_C0007099
C0007099|T047|ca in-situ|intraductal cancer_C0007099
C0007099|T047|in-situ adenocarcinoma|intraductal cancer_C0007099
C0007099|T047|in-situ ca|intraductal cancer_C0007099
C0007099|T047|in situ adenocarc|intraductal cancer_C0007099
C0007099|T047|adenoca in situ|intraductal cancer_C0007099
C0007099|T047|intraductl carc|intraductal cancer_C0007099
C0007099|T047|intraductal ca|intraductal cancer_C0007099
C0007099|T047|adenocarcinoma in situ|intraductal cancer_C0007099
C0007099|T047|adenocarcinoma in-situ|intraductal cancer_C0007099
C0007099|T047|adenocarcinoma intraductal|intraductal cancer_C0007099
C0007099|T047|adenocarcinoma intraductl|intraductal cancer_C0007099
C0007099|T047|ca intraductal|intraductal cancer_C0007099
C0007099|T047|adenoca in-situ|intraductal cancer_C0007099
C0007099|T047|intraductl cancer|intraductal cancer_C0007099
C0007099|T047|intraductl carcinoma|intraductal cancer_C0007099
C0007099|T047|adenocarc in-situ|intraductal cancer_C0007099
C0007099|T047|in-situ cancer|intraductal cancer_C0007099
C0007099|T047|intraductl adenocarcinoma|intraductal cancer_C0007099
C0007099|T047|in situ adenocarcinoma|intraductal cancer_C0007099
C0007099|T047|adenoca intraductl|intraductal cancer_C0007099
C0007099|T047|adenocarc intraductl|intraductal cancer_C0007099
C0007099|T047|adenoca intraductal|intraductal cancer_C0007099
C0007099|T047|ca in situ|intraductal cancer_C0007099
C0007099|T047|intraductl ca|intraductal cancer_C0007099
C0007099|T047|adenocarc intraductal|intraductal cancer_C0007099
C0007099|T047|in-situ carc|intraductal cancer_C0007099
C0007124|T047|in situ adenocarcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular ca in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular ca in-situ|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarc ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarc lobular|breast cancer intraductal_C0007124
C0007124|T047|lobular ca intraductl|breast cancer intraductal_C0007124
C0007124|T047|in situ ca br|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarcinoma br|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|lobular ca intraductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl cancer lobular|breast cancer intraductal_C0007124
C0007124|T047|in situ carcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|in situ ca dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarc lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarc ductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarc dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarc breast|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarc br|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenoca lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenoca ductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenoca dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenoca breast|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenoca br|breast cancer intraductal_C0007124
C0007124|T047|in situ carcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|in situ ca breast|breast cancer intraductal_C0007124
C0007124|T047|in situ carcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ carcinoma br|breast cancer intraductal_C0007124
C0007124|T047|in situ carc lobular|breast cancer intraductal_C0007124
C0007124|T047|in situ carc ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ carc dctl|breast cancer intraductal_C0007124
C0007124|T047|in situ carc breast|breast cancer intraductal_C0007124
C0007124|T047|in situ carc br|breast cancer intraductal_C0007124
C0007124|T047|in situ cancer lobular|breast cancer intraductal_C0007124
C0007124|T047|in situ cancer ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ cancer dctl|breast cancer intraductal_C0007124
C0007124|T047|in situ cancer breast|breast cancer intraductal_C0007124
C0007124|T047|in situ cancer br|breast cancer intraductal_C0007124
C0007124|T047|in situ ca lobular|breast cancer intraductal_C0007124
C0007124|T047|in situ ca ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ carcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarc dctl|breast cancer intraductal_C0007124
C0007124|T047|ductal carcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarc br|breast cancer intraductal_C0007124
C0007124|T047|dctl carc in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl carc in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl carc intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl carc intraductl|breast cancer intraductal_C0007124
C0007124|T047|dctl carcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl carcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl carcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl carcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|ductal adenoca in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal adenoca in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal adenoca intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal adenoca intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarc in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarc in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl cancer intraductl|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarc intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl cancer intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl cancer in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenoca in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenoca intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl adenoca intraductl|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarc in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarc in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarc intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarc intraductl|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl adenocarcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|dctl ca in situ|breast cancer intraductal_C0007124
C0007124|T047|dctl ca in-situ|breast cancer intraductal_C0007124
C0007124|T047|dctl ca intraductal|breast cancer intraductal_C0007124
C0007124|T047|dctl ca intraductl|breast cancer intraductal_C0007124
C0007124|T047|dctl cancer in-situ|breast cancer intraductal_C0007124
C0007124|T047|in situ adenocarc breast|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarc intraductl|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular cancer in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal carc in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal carc in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal carc intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal carc intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular cancer in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal carcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarcinoma br|breast cancer intraductal_C0007124
C0007124|T047|ductal carcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal carcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|in situ adenoca br|breast cancer intraductal_C0007124
C0007124|T047|in situ adenoca breast|breast cancer intraductal_C0007124
C0007124|T047|in situ adenoca dctl|breast cancer intraductal_C0007124
C0007124|T047|in situ adenoca ductal|breast cancer intraductal_C0007124
C0007124|T047|in situ adenoca lobular|breast cancer intraductal_C0007124
C0007124|T047|lobular cancer intraductal|breast cancer intraductal_C0007124
C0007124|T047|lobular carcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|lobular cancer intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carc in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal adenocarcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal ca in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal ca in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal ca intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal ca intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal cancer in situ|breast cancer intraductal_C0007124
C0007124|T047|ductal cancer in-situ|breast cancer intraductal_C0007124
C0007124|T047|ductal cancer intraductal|breast cancer intraductal_C0007124
C0007124|T047|ductal cancer intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carc intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular carc intraductal|breast cancer intraductal_C0007124
C0007124|T047|lobular carc in situ|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|in-situ ca dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl carcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|br ca intraductl|breast cancer intraductal_C0007124
C0007124|T047|br ca intraductal|breast cancer intraductal_C0007124
C0007124|T047|br ca in-situ|breast cancer intraductal_C0007124
C0007124|T047|br ca in situ|breast cancer intraductal_C0007124
C0007124|T047|intraductl carcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|br adenocarcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|br adenocarcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|br adenocarcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|br adenocarcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|intraductl carcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|br adenocarc intraductl|breast cancer intraductal_C0007124
C0007124|T047|br adenocarc intraductal|breast cancer intraductal_C0007124
C0007124|T047|br adenocarc in-situ|breast cancer intraductal_C0007124
C0007124|T047|br adenocarc in situ|breast cancer intraductal_C0007124
C0007124|T047|br cancer in situ|breast cancer intraductal_C0007124
C0007124|T047|br cancer in-situ|breast cancer intraductal_C0007124
C0007124|T047|br cancer intraductal|breast cancer intraductal_C0007124
C0007124|T047|br cancer intraductl|breast cancer intraductal_C0007124
C0007124|T047|intraductal cancer lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal carc br|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal carc dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal carc ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal carc lobular|breast cancer intraductal_C0007124
C0007124|T047|br carcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|intraductl carcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|br carcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|br carcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenoca in-situ|breast cancer intraductal_C0007124
C0007124|T047|br carc intraductl|breast cancer intraductal_C0007124
C0007124|T047|br carc intraductal|breast cancer intraductal_C0007124
C0007124|T047|br carc in-situ|breast cancer intraductal_C0007124
C0007124|T047|br carc in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenoca in situ|breast cancer intraductal_C0007124
C0007124|T047|br carcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|br adenoca intraductl|breast cancer intraductal_C0007124
C0007124|T047|br adenoca intraductal|breast cancer intraductal_C0007124
C0007124|T047|br adenoca in-situ|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductl ca br|breast cancer intraductal_C0007124
C0007124|T047|intraductl ca breast|breast cancer intraductal_C0007124
C0007124|T047|intraductl ca dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl ca ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl ca lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl cancer br|breast cancer intraductal_C0007124
C0007124|T047|intraductl carc ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl carc dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl carc breast|breast cancer intraductal_C0007124
C0007124|T047|intraductl carc br|breast cancer intraductal_C0007124
C0007124|T047|intraductl cancer breast|breast cancer intraductal_C0007124
C0007124|T047|intraductl cancer dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl cancer ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl carc lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal cancer ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarc lobular|breast cancer intraductal_C0007124
C0007124|T047|br adenoca in situ|breast cancer intraductal_C0007124
C0007124|T047|intraductl carcinoma br|breast cancer intraductal_C0007124
C0007124|T047|intraductal carcinoma br|breast cancer intraductal_C0007124
C0007124|T047|intraductal carcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal carcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal carcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal carcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarcinoma br|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenoca br|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenoca dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenoca ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenoca lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarc br|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarc breast|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarc dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenocarc ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductl adenoca breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal cancer dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal carc breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal cancer br|breast cancer intraductal_C0007124
C0007124|T047|breast carcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast carcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast carcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast carcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarcinoma in situ|breast cancer intraductal_C0007124
C0007124|T047|breast carc intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast carc intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast carc in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast carc in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarc intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast cancer intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast cancer intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast cancer in-situ|breast cancer intraductal_C0007124
C0007124|T047|intraductal cancer breast|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarc intraductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ carcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ carcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ carcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ carcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|in-situ adenocarcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ ca br|breast cancer intraductal_C0007124
C0007124|T047|in-situ ca breast|breast cancer intraductal_C0007124
C0007124|T047|in-situ ca ductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ ca lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ cancer br|breast cancer intraductal_C0007124
C0007124|T047|in-situ cancer breast|breast cancer intraductal_C0007124
C0007124|T047|breast ca intraductl|breast cancer intraductal_C0007124
C0007124|T047|in-situ cancer dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ cancer lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ carc br|breast cancer intraductal_C0007124
C0007124|T047|in-situ carc breast|breast cancer intraductal_C0007124
C0007124|T047|in-situ carc dctl|breast cancer intraductal_C0007124
C0007124|T047|in-situ carc ductal|breast cancer intraductal_C0007124
C0007124|T047|in-situ carc lobular|breast cancer intraductal_C0007124
C0007124|T047|in-situ carcinoma br|breast cancer intraductal_C0007124
C0007124|T047|in-situ cancer ductal|breast cancer intraductal_C0007124
C0007124|T047|dctl adenoca in situ|breast cancer intraductal_C0007124
C0007124|T047|breast cancer in situ|breast cancer intraductal_C0007124
C0007124|T047|breast ca in situ|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenoca br|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenoca breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenoca dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenoca ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenoca lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarc br|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarc breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarc dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarc ductal|breast cancer intraductal_C0007124
C0007124|T047|lobular adenoca intraductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarc lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarcinoma breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarcinoma dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarcinoma ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarcinoma lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal ca br|breast cancer intraductal_C0007124
C0007124|T047|intraductal ca breast|breast cancer intraductal_C0007124
C0007124|T047|intraductal ca dctl|breast cancer intraductal_C0007124
C0007124|T047|intraductal ca ductal|breast cancer intraductal_C0007124
C0007124|T047|intraductal ca lobular|breast cancer intraductal_C0007124
C0007124|T047|intraductal adenocarcinoma br|breast cancer intraductal_C0007124
C0007124|T047|breast adenoca in situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenoca in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast ca intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast adenoca intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast adenoca intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular adenoca intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarc in situ|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarc in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarc in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarc intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarc intraductl|breast cancer intraductal_C0007124
C0007124|T047|lobular adenocarc in situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarcinoma intraductl|breast cancer intraductal_C0007124
C0007124|T047|breast ca in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarcinoma intraductal|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarcinoma in-situ|breast cancer intraductal_C0007124
C0007124|T047|breast adenocarcinoma in situ|breast cancer intraductal_C0007124
C0015726|T041|Concern about Recurrence|Concern about Recurrence_C0015726
C0015726|T041|Fear of Recurrence|Concern about Recurrence_C0015726
C0024881|T061|Mastectomy|Mastectomy_C0024881
C0027627|T047|mediastatic|metastatic_C0027627
C0027627|T047|metastases|metastatic_C0027627
C0027627|T047|metastasis|metastatic_C0027627
C0027627|T047|met|metastatic_C0027627
C0027627|T047|metastatic|metastatic_C0027627
C0027627|T047|metastasize|metastatic_C0027627
C0027627|T047|matastases|metastatic_C0027627
C0027628|T047|mediastatic to lung|spread to lung_C0027628
C0027628|T047|met to lung|spread to lung_C0027628
C0027628|T047|disseminated to lung|spread to lung_C0027628
C0027628|T047|metastases to lung|spread to lung_C0027628
C0027628|T047|spread to lung|spread to lung_C0027628
C0027628|T047|metastasis to lung|spread to lung_C0027628
C0027628|T047|metastasize to lung|spread to lung_C0027628
C0027628|T047|metastatic to lung|spread to lung_C0027628
C0027629|T047|met to spine|spread to spine_C0027629
C0027629|T047|metastases to spine|spread to spine_C0027629
C0027629|T047|mediastatic to spine|spread to spine_C0027629
C0027629|T047|metastasize to spine|spread to spine_C0027629
C0027629|T047|evidence of metastatic|spread to spine_C0027629
C0027629|T047|metastasis to spine|spread to spine_C0027629
C0027629|T047|evidence of metastasis|spread to spine_C0027629
C0027629|T047|disseminated to spine|spread to spine_C0027629
C0027629|T047|evidence of metastases|spread to spine_C0027629
C0027629|T047|evidence of met|spread to spine_C0027629
C0027629|T047|evidence of mediastatic|spread to spine_C0027629
C0027629|T047|evidence of disseminated|spread to spine_C0027629
C0027629|T047|spread to spine|spread to spine_C0027629
C0027629|T047|evidence of metastasize|spread to spine_C0027629
C0027637|T047|consistent with brca|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast adenoca|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast adenocarc|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast adenocarcinoma|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast ca|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast cancer|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast carcinoma|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast origin|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast primary|consistent with metastatic breast_C0027637
C0027637|T047|consistent with metastatic|consistent with metastatic breast_C0027637
C0027637|T047|consistent with metastatic breast|consistent with metastatic breast_C0027637
C0027637|T047|consistent with breast carc|consistent with metastatic breast_C0027637
C0034804|T192|ER|ER_C0034804
C0034833|T192|PR|PR_C0034833
C0034897|T047|reoccuring|recurrent_C0034897
C0034897|T047|regional recurrence|recurrent_C0034897
C0034897|T047|recurrnet|recurrent_C0034897
C0034897|T047|recurred|recurrent_C0034897
C0034897|T047|recured|recurrent_C0034897
C0034897|T047|re currnet|recurrent_C0034897
C0034897|T047|evidence of recurrence|recurrent_C0034897
C0034897|T047|recurrent|recurrent_C0034897
C0034897|T047|recur|recurrent_C0034897
C0034897|T047|recurring|recurrent_C0034897
C0034897|T047|evidence of recur|recurrent_C0034897
C0034897|T047|recurrence|recurrent_C0034897
C0034897|T047|recuring|recurrent_C0034897
C0034897|T047|evidence of recurrent|recurrent_C0034897
C0034897|T047|local recurrence|recurrent_C0034897
C0069515|T192|HER-2|HER-2_C0069515
C0069515|T192|HER2|HER-2_C0069515
C0153690|T047|met bone|spread bony_C0153690
C0153690|T047|disseminated bone|spread bony_C0153690
C0153690|T047|spread bony|spread bony_C0153690
C0153690|T047|disseminated bony|spread bony_C0153690
C0153690|T047|bone mediastatic|spread bony_C0153690
C0153690|T047|spread bone|spread bony_C0153690
C0153690|T047|multiple bone metastasis|spread bony_C0153690
C0153690|T047|metastatic bony|spread bony_C0153690
C0153690|T047|multiple bone met|spread bony_C0153690
C0153690|T047|metastatic bone|spread bony_C0153690
C0153690|T047|metastasize bony|spread bony_C0153690
C0153690|T047|metastasize bone|spread bony_C0153690
C0153690|T047|mediastatic bone|spread bony_C0153690
C0153690|T047|metastasis bony|spread bony_C0153690
C0153690|T047|mediastatic bony|spread bony_C0153690
C0153690|T047|metastases bony|spread bony_C0153690
C0153690|T047|metastases bone|spread bony_C0153690
C0153690|T047|met bony|spread bony_C0153690
C0153690|T047|multiple bone metastases|spread bony_C0153690
C0153690|T047|bone disseminated|spread bony_C0153690
C0153690|T047|metastasis bone|spread bony_C0153690
C0153690|T047|bony mediastatic|spread bony_C0153690
C0153690|T047|bone met|spread bony_C0153690
C0153690|T047|bone mets|spread bony_C0153690
C0153690|T047|bone metastases|spread bony_C0153690
C0153690|T047|bony spread|spread bony_C0153690
C0153690|T047|bony metastatic|spread bony_C0153690
C0153690|T047|bony metastasize|spread bony_C0153690
C0153690|T047|bone metastasis|spread bony_C0153690
C0153690|T047|bony metastasis|spread bony_C0153690
C0153690|T047|bone metastatic|spread bony_C0153690
C0153690|T047|bone metastasize|spread bony_C0153690
C0153690|T047|bony metastases|spread bony_C0153690
C0153690|T047|bony mets|spread bony_C0153690
C0153690|T047|bony met|spread bony_C0153690
C0153690|T047|bony disseminated|spread bony_C0153690
C0153690|T047|bone spread|spread bony_C0153690
C0205281|T047|invasive|invasive_C0205281
C0205281|T047|infltrtng|invasive_C0205281
C0205281|T047|infiltrduct|invasive_C0205281
C0205281|T047|infiltr|invasive_C0205281
C0205281|T047|infitrating|invasive_C0205281
C0205281|T047|infil|invasive_C0205281
C0205281|T047|infiltrating|invasive_C0205281
C0206710|T191|Basal Tumor|Basal Tumor_C0206710
C0230108|T029|Infraclavicular|Infraclavicular_C0230108
C0278488|T047|br adenocarcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc disseminated|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc met|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc metastases|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc metastasis|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl spread|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal met|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal spread|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc metastasize|metastatic breast cancer_C0278488
C0278488|T047|br adenoca spread|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc spread|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal spread|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|carcinoma ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|br adenocarc metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast metastases|metastatic breast cancer_C0278488
C0278488|T047|br adenoca metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl ca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl ca disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma met|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc spread|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc met|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenocarc disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca spread|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl met|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca met|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl adenoca disseminated|metastatic breast cancer_C0278488
C0278488|T047|br adenoca metastases|metastatic breast cancer_C0278488
C0278488|T047|br adenoca metastasis|metastatic breast cancer_C0278488
C0278488|T047|br adenoca metastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast spread|metastatic breast cancer_C0278488
C0278488|T047|carc br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carc br met|metastatic breast cancer_C0278488
C0278488|T047|carc br metastases|metastatic breast cancer_C0278488
C0278488|T047|carc br metastasis|metastatic breast cancer_C0278488
C0278488|T047|carc br metastasize|metastatic breast cancer_C0278488
C0278488|T047|carc br metastatic|metastatic breast cancer_C0278488
C0278488|T047|carc br disseminated|metastatic breast cancer_C0278488
C0278488|T047|carc br spread|metastatic breast cancer_C0278488
C0278488|T047|carc breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carc breast met|metastatic breast cancer_C0278488
C0278488|T047|carc breast metastases|metastatic breast cancer_C0278488
C0278488|T047|carc breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|carc breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal spread|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl met|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl spread|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal met|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal met|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|cancer ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma met|metastatic breast cancer_C0278488
C0278488|T047|carc breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br met|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br metastases|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br metastasis|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br metastasize|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br metastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br disseminated|metastatic breast cancer_C0278488
C0278488|T047|carcinoma br spread|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast met|metastatic breast cancer_C0278488
C0278488|T047|dctl ca met|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|carcinoma breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|carc ductal spread|metastatic breast cancer_C0278488
C0278488|T047|carc ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|carc ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|carc breast spread|metastatic breast cancer_C0278488
C0278488|T047|carc dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|carc dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carc dctl met|metastatic breast cancer_C0278488
C0278488|T047|carc dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|carc dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carc dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|carc dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|carc dctl spread|metastatic breast cancer_C0278488
C0278488|T047|carc ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|carc ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|carc ductal met|metastatic breast cancer_C0278488
C0278488|T047|carc ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|carc ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|carc breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl ca metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer metastasis|metastatic breast cancer_C0278488
C0278488|T047|br adenoca met|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|disseminated breastca|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl ca|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal ca|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular ca|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic lobular carcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast tumor|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast malig|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast ca|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met dctl ca|metastatic breast cancer_C0278488
C0278488|T047|met dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|met dctl carc|metastatic breast cancer_C0278488
C0278488|T047|met dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|met ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|met ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|met ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met ductal ca|metastatic breast cancer_C0278488
C0278488|T047|met ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|met ductal carc|metastatic breast cancer_C0278488
C0278488|T047|met ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|met lobular adenoca|metastatic breast cancer_C0278488
C0278488|T047|met lobular adenocarc|metastatic breast cancer_C0278488
C0278488|T047|met lobular adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met lobular ca|metastatic breast cancer_C0278488
C0278488|T047|met lobular cancer|metastatic breast cancer_C0278488
C0278488|T047|met lobular carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastatic br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic br carc|metastatic breast cancer_C0278488
C0278488|T047|metastatic br cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic br ca|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastatic br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic br adenoca|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl ca|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl carc|metastatic breast cancer_C0278488
C0278488|T047|met lobular carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastatic br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|dctl ca metastasis|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast ca|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|dctl malig disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|br adenoca disseminated|metastatic breast cancer_C0278488
C0278488|T047|br adenoca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma met|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl carc spread|metastatic breast cancer_C0278488
C0278488|T047|dctl carc metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carc metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl malig mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carc metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl carc met|metastatic breast cancer_C0278488
C0278488|T047|dctl carc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl carc disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer spread|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer metastasize|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer met|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl cancer disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl ca spread|metastatic breast cancer_C0278488
C0278488|T047|dctl ca metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl ca metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl carc metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl malig met|metastatic breast cancer_C0278488
C0278488|T047|dctl malig metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl malig metastasis|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|disseminated brca|metastatic breast cancer_C0278488
C0278488|T047|disseminated br tumor|metastatic breast cancer_C0278488
C0278488|T047|disseminated br malignancy|metastatic breast cancer_C0278488
C0278488|T047|disseminated br malig|metastatic breast cancer_C0278488
C0278488|T047|disseminated br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated br carc|metastatic breast cancer_C0278488
C0278488|T047|disseminated br cancer|metastatic breast cancer_C0278488
C0278488|T047|disseminated br ca|metastatic breast cancer_C0278488
C0278488|T047|disseminated br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|disseminated br adenoca|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor spread|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor metastasis|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl malig metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl malig metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl malig spread|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy met|metastatic breast cancer_C0278488
C0278488|T047|disseminated breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy metastases|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy metastasize|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy metastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy spread|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor disseminated|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor mediastatic|metastatic breast cancer_C0278488
C0278488|T047|dctl tumor met|metastatic breast cancer_C0278488
C0278488|T047|dctl malignancy metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|cancer breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl spread|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|breast ca disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast ca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc spread|metastatic breast cancer_C0278488
C0278488|T047|br ca metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca metastases|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca spread|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc met|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc metastases|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc ductal spread|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast adenocarc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br ca metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast ca met|metastatic breast cancer_C0278488
C0278488|T047|breast ca metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast cancer disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast cancer mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast cancer met|metastatic breast cancer_C0278488
C0278488|T047|breast cancer metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br spread|metastatic breast cancer_C0278488
C0278488|T047|breast cancer metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast ca metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast ca metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast ca metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast ca spread|metastatic breast cancer_C0278488
C0278488|T047|br ca metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast spread|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenocarc breast spread|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca met|metastatic breast cancer_C0278488
C0278488|T047|breast adenoca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|brca spread|metastatic breast cancer_C0278488
C0278488|T047|br carc met|metastatic breast cancer_C0278488
C0278488|T047|br carc metastases|metastatic breast cancer_C0278488
C0278488|T047|br carc metastasis|metastatic breast cancer_C0278488
C0278488|T047|br carc metastasize|metastatic breast cancer_C0278488
C0278488|T047|br carc metastatic|metastatic breast cancer_C0278488
C0278488|T047|br carc spread|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br disseminated|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma met|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|br carcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast met|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br spread|metastatic breast cancer_C0278488
C0278488|T047|br cancer metastases|metastatic breast cancer_C0278488
C0278488|T047|br cancer metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br met|metastatic breast cancer_C0278488
C0278488|T047|br cancer metastasize|metastatic breast cancer_C0278488
C0278488|T047|br cancer spread|metastatic breast cancer_C0278488
C0278488|T047|br carc disseminated|metastatic breast cancer_C0278488
C0278488|T047|br carc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma br metastasis|metastatic breast cancer_C0278488
C0278488|T047|br cancer metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|br malig disseminated|metastatic breast cancer_C0278488
C0278488|T047|br malig mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br tumor mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br tumor met|metastatic breast cancer_C0278488
C0278488|T047|br tumor metastases|metastatic breast cancer_C0278488
C0278488|T047|br tumor metastasis|metastatic breast cancer_C0278488
C0278488|T047|br tumor metastasize|metastatic breast cancer_C0278488
C0278488|T047|br tumor metastatic|metastatic breast cancer_C0278488
C0278488|T047|br tumor disseminated|metastatic breast cancer_C0278488
C0278488|T047|br tumor spread|metastatic breast cancer_C0278488
C0278488|T047|brca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|brca met|metastatic breast cancer_C0278488
C0278488|T047|brca metastases|metastatic breast cancer_C0278488
C0278488|T047|brca metastasis|metastatic breast cancer_C0278488
C0278488|T047|brca metastasize|metastatic breast cancer_C0278488
C0278488|T047|brca metastatic|metastatic breast cancer_C0278488
C0278488|T047|brca disseminated|metastatic breast cancer_C0278488
C0278488|T047|br malignancy spread|metastatic breast cancer_C0278488
C0278488|T047|br malignancy metastatic|metastatic breast cancer_C0278488
C0278488|T047|br malignancy metastasize|metastatic breast cancer_C0278488
C0278488|T047|br cancer met|metastatic breast cancer_C0278488
C0278488|T047|br cancer mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br cancer disseminated|metastatic breast cancer_C0278488
C0278488|T047|br ca spread|metastatic breast cancer_C0278488
C0278488|T047|br malig met|metastatic breast cancer_C0278488
C0278488|T047|br malig metastases|metastatic breast cancer_C0278488
C0278488|T047|br malig metastasis|metastatic breast cancer_C0278488
C0278488|T047|br malig metastasize|metastatic breast cancer_C0278488
C0278488|T047|br malig metastatic|metastatic breast cancer_C0278488
C0278488|T047|br malig spread|metastatic breast cancer_C0278488
C0278488|T047|br malignancy disseminated|metastatic breast cancer_C0278488
C0278488|T047|br malignancy mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br malignancy met|metastatic breast cancer_C0278488
C0278488|T047|br malignancy metastases|metastatic breast cancer_C0278488
C0278488|T047|br malignancy metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast cancer metastasize|metastatic breast cancer_C0278488
C0278488|T047|cancer breast spread|metastatic breast cancer_C0278488
C0278488|T047|breast cancer metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast carc disseminated|metastatic breast cancer_C0278488
C0278488|T047|ca dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl spread|metastatic breast cancer_C0278488
C0278488|T047|ca dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|ca dctl spread|metastatic breast cancer_C0278488
C0278488|T047|ca ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|ca ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|ca ductal met|metastatic breast cancer_C0278488
C0278488|T047|ca ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl spread|metastatic breast cancer_C0278488
C0278488|T047|met dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|ca ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|ca breast metastases|metastatic breast cancer_C0278488
C0278488|T047|ca breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|ca breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal spread|metastatic breast cancer_C0278488
C0278488|T047|ca breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|ca breast spread|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal met|metastatic breast cancer_C0278488
C0278488|T047|ca dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|ca dctl met|metastatic breast cancer_C0278488
C0278488|T047|ca dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|ca dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|ca dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ca breast met|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl met|metastatic breast cancer_C0278488
C0278488|T047|cancer br metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer br metastasize|metastatic breast cancer_C0278488
C0278488|T047|cancer br metastatic|metastatic breast cancer_C0278488
C0278488|T047|cancer br spread|metastatic breast cancer_C0278488
C0278488|T047|cancer breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|cancer breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca br spread|metastatic breast cancer_C0278488
C0278488|T047|cancer breast met|metastatic breast cancer_C0278488
C0278488|T047|adenoca br metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca br metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenoca br metastases|metastatic breast cancer_C0278488
C0278488|T047|cancer breast metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|cancer breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca br metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast met|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast spread|metastatic breast cancer_C0278488
C0278488|T047|ca ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|ca ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|ca ductal spread|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|cancer br disseminated|metastatic breast cancer_C0278488
C0278488|T047|cancer br met|metastatic breast cancer_C0278488
C0278488|T047|cancer br metastases|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenoca breast metastases|metastatic breast cancer_C0278488
C0278488|T047|cancer br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ca breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ca breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|ca br spread|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma met|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast carc spread|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast malig disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast malig mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast malig met|metastatic breast cancer_C0278488
C0278488|T047|breast malig metastases|metastatic breast cancer_C0278488
C0278488|T047|breast malig metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast malig metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast carcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|breast malig metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast carc metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast carc metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast carc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarcinoma dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|br ca metastases|metastatic breast cancer_C0278488
C0278488|T047|br ca met|metastatic breast cancer_C0278488
C0278488|T047|br ca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast carc met|metastatic breast cancer_C0278488
C0278488|T047|breast carc metastasize|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br metastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br metastasis|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br met|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast carc metastases|metastatic breast cancer_C0278488
C0278488|T047|adenocarc br metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast malig spread|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|breastca met|metastatic breast cancer_C0278488
C0278488|T047|breastca metastases|metastatic breast cancer_C0278488
C0278488|T047|breastca metastasis|metastatic breast cancer_C0278488
C0278488|T047|breastca metastasize|metastatic breast cancer_C0278488
C0278488|T047|breastca metastatic|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|breastca spread|metastatic breast cancer_C0278488
C0278488|T047|ca br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ca br met|metastatic breast cancer_C0278488
C0278488|T047|ca br metastases|metastatic breast cancer_C0278488
C0278488|T047|ca br metastasis|metastatic breast cancer_C0278488
C0278488|T047|ca br metastasize|metastatic breast cancer_C0278488
C0278488|T047|ca br metastatic|metastatic breast cancer_C0278488
C0278488|T047|ca br disseminated|metastatic breast cancer_C0278488
C0278488|T047|breastca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|br adenocarcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|br ca disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy met|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy metastases|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast malignancy spread|metastatic breast cancer_C0278488
C0278488|T047|breast tumor disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast tumor mediastatic|metastatic breast cancer_C0278488
C0278488|T047|breast tumor met|metastatic breast cancer_C0278488
C0278488|T047|breast tumor metastases|metastatic breast cancer_C0278488
C0278488|T047|breast tumor metastasis|metastatic breast cancer_C0278488
C0278488|T047|breast tumor metastasize|metastatic breast cancer_C0278488
C0278488|T047|breast tumor metastatic|metastatic breast cancer_C0278488
C0278488|T047|breast tumor spread|metastatic breast cancer_C0278488
C0278488|T047|breastca disseminated|metastatic breast cancer_C0278488
C0278488|T047|breast cancer spread|metastatic breast cancer_C0278488
C0278488|T047|met dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis br adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasis breastca|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast malig|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast carc|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast ca|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasis breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasis brca|metastatic breast cancer_C0278488
C0278488|T047|metastasis br tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasis br malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasis br malig|metastatic breast cancer_C0278488
C0278488|T047|metastasis br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis br carc|metastatic breast cancer_C0278488
C0278488|T047|metastasis br cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasis br ca|metastatic breast cancer_C0278488
C0278488|T047|metastasis br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|met dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl ca|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize brca|metastatic breast cancer_C0278488
C0278488|T047|metastasize br tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasize br malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasize br malig|metastatic breast cancer_C0278488
C0278488|T047|metastasize br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize br carc|metastatic breast cancer_C0278488
C0278488|T047|metastasize br cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize br ca|metastatic breast cancer_C0278488
C0278488|T047|metastasize br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasize br adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal malig|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal carc|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal ca|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl malig|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasis dctl carc|metastatic breast cancer_C0278488
C0278488|T047|metastasis ductal malig|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|metastases br carc|metastatic breast cancer_C0278488
C0278488|T047|metastases br cancer|metastatic breast cancer_C0278488
C0278488|T047|metastases br ca|metastatic breast cancer_C0278488
C0278488|T047|metastases br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastases br adenoca|metastatic breast cancer_C0278488
C0278488|T047|met ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|met ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|met ductal malig|metastatic breast cancer_C0278488
C0278488|T047|met dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|met dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|met dctl malig|metastatic breast cancer_C0278488
C0278488|T047|met breastca|metastatic breast cancer_C0278488
C0278488|T047|met breast tumor|metastatic breast cancer_C0278488
C0278488|T047|met breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|met breast malig|metastatic breast cancer_C0278488
C0278488|T047|met brca|metastatic breast cancer_C0278488
C0278488|T047|met br tumor|metastatic breast cancer_C0278488
C0278488|T047|met br malignancy|metastatic breast cancer_C0278488
C0278488|T047|met br malig|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular carc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases br malig|metastatic breast cancer_C0278488
C0278488|T047|metastases br malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastases br tumor|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal ca|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl malig|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl carc|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl ca|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases ductal carc|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastases breastca|metastatic breast cancer_C0278488
C0278488|T047|metastases breast tumor|metastatic breast cancer_C0278488
C0278488|T047|metastases breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastases breast malig|metastatic breast cancer_C0278488
C0278488|T047|metastases breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases breast carc|metastatic breast cancer_C0278488
C0278488|T047|metastases breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastases breast ca|metastatic breast cancer_C0278488
C0278488|T047|metastases breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastases breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastases breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastases brca|metastatic breast cancer_C0278488
C0278488|T047|metastases dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast ca|metastatic breast cancer_C0278488
C0278488|T047|tumor br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor br disseminated|metastatic breast cancer_C0278488
C0278488|T047|spread ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|spread ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|spread ductal malig|metastatic breast cancer_C0278488
C0278488|T047|spread ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread ductal carc|metastatic breast cancer_C0278488
C0278488|T047|spread ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|spread ductal ca|metastatic breast cancer_C0278488
C0278488|T047|spread ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|spread ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|spread dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|spread dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|spread dctl malig|metastatic breast cancer_C0278488
C0278488|T047|spread dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread dctl carc|metastatic breast cancer_C0278488
C0278488|T047|spread dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|spread dctl ca|metastatic breast cancer_C0278488
C0278488|T047|spread dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|spread dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|spread breastca|metastatic breast cancer_C0278488
C0278488|T047|spread breast tumor|metastatic breast cancer_C0278488
C0278488|T047|spread breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|tumor br met|metastatic breast cancer_C0278488
C0278488|T047|tumor br metastases|metastatic breast cancer_C0278488
C0278488|T047|tumor br metastasis|metastatic breast cancer_C0278488
C0278488|T047|tumor br metastasize|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal spread|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal met|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl spread|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|spread breast malig|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|tumor breast spread|metastatic breast cancer_C0278488
C0278488|T047|tumor breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|tumor breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|tumor breast metastases|metastatic breast cancer_C0278488
C0278488|T047|tumor breast met|metastatic breast cancer_C0278488
C0278488|T047|tumor breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|tumor br spread|metastatic breast cancer_C0278488
C0278488|T047|tumor br metastatic|metastatic breast cancer_C0278488
C0278488|T047|tumor dctl met|metastatic breast cancer_C0278488
C0278488|T047|spread breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread breast carc|metastatic breast cancer_C0278488
C0278488|T047|spread breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal malig|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal carc|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal ca|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl malig|metastatic breast cancer_C0278488
C0278488|T047|metastasize ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl ca|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastasize breastca|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast tumor|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast malig|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast carc|metastatic breast cancer_C0278488
C0278488|T047|metastasize breast cancer|metastatic breast cancer_C0278488
C0278488|T047|metastasize dctl carc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular adenocarc|metastatic breast cancer_C0278488
C0278488|T047|metastatic br malig|metastatic breast cancer_C0278488
C0278488|T047|metastatic br tumor|metastatic breast cancer_C0278488
C0278488|T047|spread breast ca|metastatic breast cancer_C0278488
C0278488|T047|spread breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|spread breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|spread brca|metastatic breast cancer_C0278488
C0278488|T047|spread br tumor|metastatic breast cancer_C0278488
C0278488|T047|spread br malignancy|metastatic breast cancer_C0278488
C0278488|T047|spread br malig|metastatic breast cancer_C0278488
C0278488|T047|spread br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread br carc|metastatic breast cancer_C0278488
C0278488|T047|spread br cancer|metastatic breast cancer_C0278488
C0278488|T047|spread br ca|metastatic breast cancer_C0278488
C0278488|T047|metastatic br malignancy|metastatic breast cancer_C0278488
C0278488|T047|spread br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|spread br adenoca|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastatic ductal malig|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastatic dctl malig|metastatic breast cancer_C0278488
C0278488|T047|metastatic breastca|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast tumor|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|metastatic breast malig|metastatic breast cancer_C0278488
C0278488|T047|metastatic brca|metastatic breast cancer_C0278488
C0278488|T047|spread br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic lobular adenoca|metastatic breast cancer_C0278488
C0278488|T047|met br adenoca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal carc|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal malig|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal malignancy|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy spread|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca met|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy met|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenoca spread|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc met|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor met|metastatic breast cancer_C0278488
C0278488|T047|malig breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|malig breast met|metastatic breast cancer_C0278488
C0278488|T047|malig breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malig breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|malig br spread|metastatic breast cancer_C0278488
C0278488|T047|malig br metastatic|metastatic breast cancer_C0278488
C0278488|T047|malig br metastasize|metastatic breast cancer_C0278488
C0278488|T047|malig br metastasis|metastatic breast cancer_C0278488
C0278488|T047|malig br metastases|metastatic breast cancer_C0278488
C0278488|T047|malig br met|metastatic breast cancer_C0278488
C0278488|T047|malig br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malig br disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor spread|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor metastasis|metastatic breast cancer_C0278488
C0278488|T047|met br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|ductal tumor metastases|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|disseminated ductal ca|metastatic breast cancer_C0278488
C0278488|T047|malig breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal malignancy disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal malig metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal carc disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer spread|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer met|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal cancer disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal ca spread|metastatic breast cancer_C0278488
C0278488|T047|ductal ca metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal ca metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal ca metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal ca metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal ca met|metastatic breast cancer_C0278488
C0278488|T047|ductal ca mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal ca disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal carc mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal malig spread|metastatic breast cancer_C0278488
C0278488|T047|ductal carc met|metastatic breast cancer_C0278488
C0278488|T047|ductal carc metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal malig metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal malig metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal malig metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal malig met|metastatic breast cancer_C0278488
C0278488|T047|ductal malig mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal malig disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma spread|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma metastasis|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma metastases|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma met|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma mediastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal carcinoma disseminated|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal carc spread|metastatic breast cancer_C0278488
C0278488|T047|ductal carc metastatic|metastatic breast cancer_C0278488
C0278488|T047|ductal carc metastasize|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal tumor|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarc spread|metastatic breast cancer_C0278488
C0278488|T047|ductal carc metastases|metastatic breast cancer_C0278488
C0278488|T047|malig breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|malig breast metastases|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast malig|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast carc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|met breast adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met breast adenocarc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic brca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast malignancy|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br tumor|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br malig|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br carc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br adenocarc|metastatic breast cancer_C0278488
C0278488|T047|met breast adenoca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br adenoca|metastatic breast cancer_C0278488
C0278488|T047|met br carcinoma|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal spread|metastatic breast cancer_C0278488
C0278488|T047|mediastatic br malignancy|metastatic breast cancer_C0278488
C0278488|T047|malig breast spread|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breast tumor|metastatic breast cancer_C0278488
C0278488|T047|met breast ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal malig|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal carc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal adenocarc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic ductal adenoca|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl malig|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|mediastatic breastca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl malignancy|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl carc|metastatic breast cancer_C0278488
C0278488|T047|disseminated dctl tumor|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl ca|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl adenocarcinoma|metastatic breast cancer_C0278488
C0278488|T047|met breast carcinoma|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl adenocarc|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl adenoca|metastatic breast cancer_C0278488
C0278488|T047|met breast carc|metastatic breast cancer_C0278488
C0278488|T047|met breast cancer|metastatic breast cancer_C0278488
C0278488|T047|mediastatic dctl malig|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|ductal adenocarcinoma met|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|malignancy br metastasize|metastatic breast cancer_C0278488
C0278488|T047|malignancy br metastasis|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|malignancy br met|metastatic breast cancer_C0278488
C0278488|T047|malignancy br mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy br disseminated|metastatic breast cancer_C0278488
C0278488|T047|malig ductal spread|metastatic breast cancer_C0278488
C0278488|T047|malig ductal metastatic|metastatic breast cancer_C0278488
C0278488|T047|malig ductal metastasize|metastatic breast cancer_C0278488
C0278488|T047|malig ductal metastasis|metastatic breast cancer_C0278488
C0278488|T047|malignancy br metastatic|metastatic breast cancer_C0278488
C0278488|T047|malig ductal metastases|metastatic breast cancer_C0278488
C0278488|T047|malig ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malig ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|malig dctl spread|metastatic breast cancer_C0278488
C0278488|T047|malig dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|malig dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|malig dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|malig dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|malig dctl met|metastatic breast cancer_C0278488
C0278488|T047|malig dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malig dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|malig ductal met|metastatic breast cancer_C0278488
C0278488|T047|malignancy br spread|metastatic breast cancer_C0278488
C0278488|T047|malignancy br metastases|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal met|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy ductal disseminated|metastatic breast cancer_C0278488
C0278488|T047|met br carc|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl spread|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl metastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl metastasize|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl metastasis|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl metastases|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl met|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast disseminated|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl disseminated|metastatic breast cancer_C0278488
C0278488|T047|malignancy dctl mediastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast metastatic|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast met|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast metastases|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast metastasis|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast spread|metastatic breast cancer_C0278488
C0278488|T047|malignancy breast metastasize|metastatic breast cancer_C0278488
C0278488|T047|met br ca|metastatic breast cancer_C0278488
C0278488|T047|met br cancer|metastatic breast cancer_C0278488
C0278489|T047|br metastatic|metastatic breast_C0278489
C0278489|T047|br met|metastatic breast_C0278489
C0278489|T047|br spread|metastatic breast_C0278489
C0278489|T047|br metastasize|metastatic breast_C0278489
C0278489|T047|br disseminated|metastatic breast_C0278489
C0278489|T047|disseminated ductal|metastatic breast_C0278489
C0278489|T047|br mediastatic|metastatic breast_C0278489
C0278489|T047|spread ductal|metastatic breast_C0278489
C0278489|T047|disseminated dctl|metastatic breast_C0278489
C0278489|T047|br metastasis|metastatic breast_C0278489
C0278489|T047|br metastases|metastatic breast_C0278489
C0278489|T047|spread br|metastatic breast_C0278489
C0278489|T047|spread breast|metastatic breast_C0278489
C0278489|T047|breast met|metastatic breast_C0278489
C0278489|T047|breast metastases|metastatic breast_C0278489
C0278489|T047|breast metastasis|metastatic breast_C0278489
C0278489|T047|breast metastasize|metastatic breast_C0278489
C0278489|T047|breast metastatic|metastatic breast_C0278489
C0278489|T047|breast spread|metastatic breast_C0278489
C0278489|T047|metastasize br|metastatic breast_C0278489
C0278489|T047|metastasis ductal|metastatic breast_C0278489
C0278489|T047|metastasis dctl|metastatic breast_C0278489
C0278489|T047|metastasis breast|metastatic breast_C0278489
C0278489|T047|metastasis br|metastatic breast_C0278489
C0278489|T047|metastases ductal|metastatic breast_C0278489
C0278489|T047|mediastatic br|metastatic breast_C0278489
C0278489|T047|metastases dctl|metastatic breast_C0278489
C0278489|T047|mediastatic breast|metastatic breast_C0278489
C0278489|T047|metastases breast|metastatic breast_C0278489
C0278489|T047|metastases br|metastatic breast_C0278489
C0278489|T047|mediastatic dctl|metastatic breast_C0278489
C0278489|T047|met ductal|metastatic breast_C0278489
C0278489|T047|met dctl|metastatic breast_C0278489
C0278489|T047|met breast|metastatic breast_C0278489
C0278489|T047|met br|metastatic breast_C0278489
C0278489|T047|spread dctl|metastatic breast_C0278489
C0278489|T047|breast mediastatic|metastatic breast_C0278489
C0278489|T047|dctl disseminated|metastatic breast_C0278489
C0278489|T047|mediastatic ductal|metastatic breast_C0278489
C0278489|T047|ductal spread|metastatic breast_C0278489
C0278489|T047|disseminated breast|metastatic breast_C0278489
C0278489|T047|metastasize breast|metastatic breast_C0278489
C0278489|T047|metastatic ductal|metastatic breast_C0278489
C0278489|T047|metastatic breast|metastatic breast_C0278489
C0278489|T047|disseminated br|metastatic breast_C0278489
C0278489|T047|ductal disseminated|metastatic breast_C0278489
C0278489|T047|metastatic br|metastatic breast_C0278489
C0278489|T047|dctl spread|metastatic breast_C0278489
C0278489|T047|dctl metastatic|metastatic breast_C0278489
C0278489|T047|metastasize ductal|metastatic breast_C0278489
C0278489|T047|dctl metastasize|metastatic breast_C0278489
C0278489|T047|dctl metastasis|metastatic breast_C0278489
C0278489|T047|metastatic dctl|metastatic breast_C0278489
C0278489|T047|dctl metastases|metastatic breast_C0278489
C0278489|T047|dctl met|metastatic breast_C0278489
C0278489|T047|dctl mediastatic|metastatic breast_C0278489
C0278489|T047|breast disseminated|metastatic breast_C0278489
C0278489|T047|ductal metastatic|metastatic breast_C0278489
C0278489|T047|metastasize dctl|metastatic breast_C0278489
C0278489|T047|ductal mediastatic|metastatic breast_C0278489
C0278489|T047|ductal met|metastatic breast_C0278489
C0278489|T047|ductal metastases|metastatic breast_C0278489
C0278489|T047|ductal metastasize|metastatic breast_C0278489
C0278489|T047|ductal metastasis|metastatic breast_C0278489
C0278493|T047|lobular recurrnet cancer|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet carc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet cancer|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet cancer|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrnet adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrnet adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet ca|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet adenoca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet cancer|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recur br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recur breast|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrnet adenoca|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet adenoca|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|br recurrnet carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrnet lobular|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrnet ductal|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrnet dctl|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrnet br|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet ca|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrnet adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrnet breast|recurrnet breast cancer_C0278493
C0278493|T047|recurrnet lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence cancer|recurrnet breast cancer_C0278493
C0278493|T047|ca recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence adenoca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring carc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring cancer|recurrnet breast cancer_C0278493
C0278493|T047|ca recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ca recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur carc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur cancer|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur ca|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ca recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|ca recurring br|recurrnet breast cancer_C0278493
C0278493|T047|ca recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|ca recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|lobular recuring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ca recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|ca recuring br|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence ca|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence adenoca|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring ca|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ca recur br|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence carc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrence carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent adenoca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ca recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|ca recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|ca recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|ca recur breast|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurrent adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrence carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring ca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast carc|recurrnet breast cancer_C0278493
C0278493|T047|ca recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recur br|recurrnet breast cancer_C0278493
C0278493|T047|cancer recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|cancer recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|cancer recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|cancer recuring br|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|breast recur carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|cancer recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recur carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recur cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recur ca|recurrnet breast cancer_C0278493
C0278493|T047|breast recur adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recur adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|cancer recur breast|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br carc|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence carc|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recuring br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurring br|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring cancer|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recur breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recur br|recurrnet breast cancer_C0278493
C0278493|T047|lobular recur adenoca|recurrnet breast cancer_C0278493
C0278493|T047|breast recuring carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|ca recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent adenoca|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring br ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast ca|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring br cancer|recurrnet breast cancer_C0278493
C0278493|T047|recuring br carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast ca|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast carc|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recuring dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recuring breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recuring br|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent carc|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent ca|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenoca recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring carc|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring cancer|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring ca|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|lobular recurring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrence lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|recurring dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurring lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur breast carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur breast carc|recurrnet breast cancer_C0278493
C0278493|T047|recur breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrence dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurring ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrence breast carc|recurrnet breast cancer_C0278493
C0278493|T047|recur br ca|recurrnet breast cancer_C0278493
C0278493|T047|recur br carc|recurrnet breast cancer_C0278493
C0278493|T047|recur br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recur breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recur breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recur breast ca|recurrnet breast cancer_C0278493
C0278493|T047|recur br cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl adenoca|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence adenoca|recurrnet breast cancer_C0278493
C0278493|T047|br recuring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recuring carc|recurrnet breast cancer_C0278493
C0278493|T047|br recuring cancer|recurrnet breast cancer_C0278493
C0278493|T047|br recuring ca|recurrnet breast cancer_C0278493
C0278493|T047|br recuring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recuring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recur carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recur carc|recurrnet breast cancer_C0278493
C0278493|T047|br recur cancer|recurrnet breast cancer_C0278493
C0278493|T047|br recur ca|recurrnet breast cancer_C0278493
C0278493|T047|br recur adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recur adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recuring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal cancer|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recurring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal ca|recurrnet breast cancer_C0278493
C0278493|T047|br recurring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recurring ca|recurrnet breast cancer_C0278493
C0278493|T047|br recurring cancer|recurrnet breast cancer_C0278493
C0278493|T047|br recurring carc|recurrnet breast cancer_C0278493
C0278493|T047|br recurring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|breast recur adenoca|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence ca|recurrnet breast cancer_C0278493
C0278493|T047|br recurring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal carc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular adenoca|recurrnet breast cancer_C0278493
C0278493|T047|carc recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|carc recuring br|recurrnet breast cancer_C0278493
C0278493|T047|carc recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|carc recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|carc recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|carc recur breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|carc recur br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular carc|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|carc recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular ca|recurrnet breast cancer_C0278493
C0278493|T047|br recur adenoca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurring br|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular cancer|recurrnet breast cancer_C0278493
C0278493|T047|breast recurrent carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast cancer|recurrnet breast cancer_C0278493
C0278493|T047|carc recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent carc|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent cancer|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recur breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recur br|recurrnet breast cancer_C0278493
C0278493|T047|carc recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recuring br|recurrnet breast cancer_C0278493
C0278493|T047|carc recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|carc recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|carc recurring br|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur ca|recurrnet breast cancer_C0278493
C0278493|T047|carc recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurring br|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|carcinoma recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur cancer|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring cancer|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring carc|recurrnet breast cancer_C0278493
C0278493|T047|carc recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|br recurrence carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent adenoca|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|br recurrent ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent cancer|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring cancer|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recuring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence ca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence cancer|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence carc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrence carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent adenoca|recurrnet breast cancer_C0278493
C0278493|T047|dctl recurrent adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|dctl recur carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurring br|recurrnet breast cancer_C0278493
C0278493|T047|carc recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recur br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recur ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recur lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recuring br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recuring breast|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurring dctl|recurrnet breast cancer_C0278493
C0278493|T047|recurring br carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recur dctl|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl carc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent adenoca|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|cancer recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring cancer|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring carc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recur breast|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring cancer|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring carc|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence cancer|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence carc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring br ca|recurrnet breast cancer_C0278493
C0278493|T047|recurring br cancer|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrent breast|recurrnet breast cancer_C0278493
C0278493|T047|recurring br carc|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrent br|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrence lobular|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurring ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrence ca|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur carc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur cancer|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur ca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent carc|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurring br|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal adenoca|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent ductal adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurring breast|recurrnet breast cancer_C0278493
C0278493|T047|recurrent lobular carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrence breast|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent cancer|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrence ductal|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurring ductal|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrent lobular|recurrnet breast cancer_C0278493
C0278493|T047|recurrent dctl carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrent ductal|recurrnet breast cancer_C0278493
C0278493|T047|recurring br adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring br adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|recurring br adenoca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurrence dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recuring dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recuring lobular|recurrnet breast cancer_C0278493
C0278493|T047|ductal recuring adenoca|recurrnet breast cancer_C0278493
C0278493|T047|ductal recurrent ca|recurrnet breast cancer_C0278493
C0278493|T047|adenocarc recurring lobular|recurrnet breast cancer_C0278493
C0278493|T047|ductal recur carcinoma|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrent dctl|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recurrence br|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast adenocarcinoma|recurrnet breast cancer_C0278493
C0278493|T047|recurring breast adenocarc|recurrnet breast cancer_C0278493
C0278493|T047|adenocarcinoma recuring ductal|recurrnet breast cancer_C0278493
C0278493|T047|cancer recurrent breast|recurrnet breast cancer_C0278493
C0278588|T047|newly diagnosed met brca|newly diagnosed metastatic breast cancer_C0278588
C0278588|T047|newly diagnosed metastatic breast cancer|newly diagnosed metastatic breast cancer_C0278588
C0278588|T047|newly diagnosed metastatic breast ca|newly diagnosed metastatic breast cancer_C0278588
C0278588|T047|newly diagnosed metastatic brca|newly diagnosed metastatic breast cancer_C0278588
C0278588|T047|newly diagnosed met breast ca|newly diagnosed metastatic breast cancer_C0278588
C0278588|T047|newly diagnosed met breast cancer|newly diagnosed metastatic breast cancer_C0278588
C0343834|T047|bone lesion|bone lesion_C0343834
C0343834|T047|bony lesion|bone lesion_C0343834
C0343834|T047|lesion bone|bone lesion_C0343834
C0343834|T047|lesion bony|bone lesion_C0343834
C0343835|T047|met lesion|metastatic lesion_C0343835
C0343835|T047|metastatic lesion|metastatic lesion_C0343835
C0438105|T047|carcinoma br reoccur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast recur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl recur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast progressive|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|recurrent breast tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrent breastca|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer progressive|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl ca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl ca reoccur|recurrent breast cancer_C0438105
C0438105|T047|recurrence br malignancy|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer recur|recurrent breast cancer_C0438105
C0438105|T047|recurrence br malig|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl ca recur|recurrent breast cancer_C0438105
C0438105|T047|dctl ca recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl ca recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl ca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl ca progressive|recurrent breast cancer_C0438105
C0438105|T047|chest wall recur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca progressive|recurrent breast cancer_C0438105
C0438105|T047|recurrent br tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccur br malig|recurrent breast cancer_C0438105
C0438105|T047|reoccur br carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur br carc|recurrent breast cancer_C0438105
C0438105|T047|reoccur br cancer|recurrent breast cancer_C0438105
C0438105|T047|reoccur br ca|recurrent breast cancer_C0438105
C0438105|T047|reoccur br adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur br adenocarc|recurrent breast cancer_C0438105
C0438105|T047|recurrent br malignancy|recurrent breast cancer_C0438105
C0438105|T047|recurrent br malig|recurrent breast cancer_C0438105
C0438105|T047|recurrence ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrence ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|recurrence ductal malig|recurrent breast cancer_C0438105
C0438105|T047|recurrence dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccur br adenoca|recurrent breast cancer_C0438105
C0438105|T047|recurrence dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|chest wall recurrence|recurrent breast cancer_C0438105
C0438105|T047|chest wall recurrent|recurrent breast cancer_C0438105
C0438105|T047|recurrent dctl malig|recurrent breast cancer_C0438105
C0438105|T047|recurrent dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|recurrence brca|recurrent breast cancer_C0438105
C0438105|T047|recurrence breast malig|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca recur|recurrent breast cancer_C0438105
C0438105|T047|recurrent dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrent ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|recurrent ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrence breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|recurrence breast tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrence breastca|recurrent breast cancer_C0438105
C0438105|T047|recurrence dctl malig|recurrent breast cancer_C0438105
C0438105|T047|recurrent ductal malig|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca recurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccur br malignancy|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc recurrent|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc recur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenocarc progressive|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br recurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br recur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal recur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|carcinoma br progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccur br tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrent brca|recurrent breast cancer_C0438105
C0438105|T047|reoccur brca|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca recurrent|recurrent breast cancer_C0438105
C0438105|T047|recurrent breast malig|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|carcinoma ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl adenoca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|recurrence br tumor|recurrent breast cancer_C0438105
C0438105|T047|recurrent breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal malig progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal malig recur|recurrent breast cancer_C0438105
C0438105|T047|ductal malig recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal malig recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal malig reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal malig reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal malig reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy recur|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal malignancy reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor recur|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal tumor reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal ca progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal ca recur|recurrent breast cancer_C0438105
C0438105|T047|ductal ca recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal ca recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal ca reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal ca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal ca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer recur|recurrent breast cancer_C0438105
C0438105|T047|malig br progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal carc progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal carc recur|recurrent breast cancer_C0438105
C0438105|T047|ductal carc recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal carc recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal carc reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal carc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal carc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal carcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal cancer recurrent|recurrent breast cancer_C0438105
C0438105|T047|malig br recur|recurrent breast cancer_C0438105
C0438105|T047|malig br recurrence|recurrent breast cancer_C0438105
C0438105|T047|malig br recurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy br reoccur|recurrent breast cancer_C0438105
C0438105|T047|malignancy br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast progressive|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast recur|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|malignancy br recurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl recur|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal recur|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malignancy dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|malignancy br recurrence|recurrent breast cancer_C0438105
C0438105|T047|malignancy br progressive|recurrent breast cancer_C0438105
C0438105|T047|malig br reoccur|recurrent breast cancer_C0438105
C0438105|T047|malig br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malig br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malig breast progressive|recurrent breast cancer_C0438105
C0438105|T047|malig breast recur|recurrent breast cancer_C0438105
C0438105|T047|malig breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|malig breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|malig breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|malig breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malig breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malig dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|malignancy br recur|recurrent breast cancer_C0438105
C0438105|T047|malig dctl recur|recurrent breast cancer_C0438105
C0438105|T047|malig dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|malig dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|malig dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malig dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malig ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|malig ductal recur|recurrent breast cancer_C0438105
C0438105|T047|malig ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|malig ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|malig ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|malig ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|malig ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|malig dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|recur ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|recur ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|recur ductal malig|recurrent breast cancer_C0438105
C0438105|T047|recur dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|recur dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|recur dctl malig|recurrent breast cancer_C0438105
C0438105|T047|recur breastca|recurrent breast cancer_C0438105
C0438105|T047|recur breast tumor|recurrent breast cancer_C0438105
C0438105|T047|recur breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy reoccur|recurrent breast cancer_C0438105
C0438105|T047|recur breast malig|recurrent breast cancer_C0438105
C0438105|T047|recur br tumor|recurrent breast cancer_C0438105
C0438105|T047|recur br malignancy|recurrent breast cancer_C0438105
C0438105|T047|recur br malig|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor recur|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl tumor reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|recur brca|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy recur|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl carc progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl carc recur|recurrent breast cancer_C0438105
C0438105|T047|dctl carc recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl carc recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl carc reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl carc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl carc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl malig progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl malig recur|recurrent breast cancer_C0438105
C0438105|T047|dctl malig recurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl malig recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl malig reoccur|recurrent breast cancer_C0438105
C0438105|T047|dctl malig reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|dctl malig reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl malignancy progressive|recurrent breast cancer_C0438105
C0438105|T047|dctl carcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|dctl cancer recurrent|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal malig|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal carc|recurrent breast cancer_C0438105
C0438105|T047|progressive br malignancy|recurrent breast cancer_C0438105
C0438105|T047|progressive br malig|recurrent breast cancer_C0438105
C0438105|T047|progressive br carcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive br carc|recurrent breast cancer_C0438105
C0438105|T047|progressive br cancer|recurrent breast cancer_C0438105
C0438105|T047|progressive br ca|recurrent breast cancer_C0438105
C0438105|T047|progressive br adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive br adenocarc|recurrent breast cancer_C0438105
C0438105|T047|progressive br adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast ca|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca recur|recurrent breast cancer_C0438105
C0438105|T047|progressive br tumor|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc recur|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc recurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc recurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc reoccur|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ductal adenocarcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|ductal adenoca recurrent|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal carcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive brca|recurrent breast cancer_C0438105
C0438105|T047|progressive breast adenocarc|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal cancer|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal ca|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal adenocarc|recurrent breast cancer_C0438105
C0438105|T047|progressive ductal adenoca|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl malig|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl carcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl carc|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl cancer|recurrent breast cancer_C0438105
C0438105|T047|progressive breast adenoca|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl ca|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl adenocarc|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl adenoca|recurrent breast cancer_C0438105
C0438105|T047|progressive breastca|recurrent breast cancer_C0438105
C0438105|T047|progressive breast tumor|recurrent breast cancer_C0438105
C0438105|T047|progressive breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|progressive breast malig|recurrent breast cancer_C0438105
C0438105|T047|progressive breast carcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive breast carc|recurrent breast cancer_C0438105
C0438105|T047|progressive breast cancer|recurrent breast cancer_C0438105
C0438105|T047|progressive breast ca|recurrent breast cancer_C0438105
C0438105|T047|progressive breast adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|progressive dctl adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast cancer|recurrent breast cancer_C0438105
C0438105|T047|carcinoma dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast carcinoma|recurrent breast cancer_C0438105
C0438105|T047|breast malig reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast malig reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast malig recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast malig recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast malig recur|recurrent breast cancer_C0438105
C0438105|T047|breast malig progressive|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast malig reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|breast carc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast carc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast carc reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast carcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast carc recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy progressive|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy recurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal ca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal cancer|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy recur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal malig|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast malignancy recurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent ductal carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl malig|recurrent breast cancer_C0438105
C0438105|T047|breast carc recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast carc progressive|recurrent breast cancer_C0438105
C0438105|T047|breast ca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast ca reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast ca recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast ca recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast ca recur|recurrent breast cancer_C0438105
C0438105|T047|breast ca progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast ca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|breast carc recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast cancer reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast cancer reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast cancer reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast cancer recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast cancer recur|recurrent breast cancer_C0438105
C0438105|T047|breast cancer progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc breast recur|recurrent breast cancer_C0438105
C0438105|T047|breast cancer recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl cancer|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal recur|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ca breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br cancer|recurrent breast cancer_C0438105
C0438105|T047|ca breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ca breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|ca breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|ca breast recur|recurrent breast cancer_C0438105
C0438105|T047|ca breast progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br carcinoma|recurrent breast cancer_C0438105
C0438105|T047|ca breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br malig|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ca dctl recur|recurrent breast cancer_C0438105
C0438105|T047|ca ductal recur|recurrent breast cancer_C0438105
C0438105|T047|ca ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl recur|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|ca dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br ca|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ca dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|ca dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ca dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|ca dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|ca dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenoca dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br malignancy|recurrent breast cancer_C0438105
C0438105|T047|ca br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast carcinoma|recurrent breast cancer_C0438105
C0438105|T047|breast tumor reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast tumor reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast tumor reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast tumor recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast tumor recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast tumor recur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast carc|recurrent breast cancer_C0438105
C0438105|T047|breast tumor progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breastca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl ca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast malig|recurrent breast cancer_C0438105
C0438105|T047|ca br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast cancer|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|ca br reoccur|recurrent breast cancer_C0438105
C0438105|T047|ca br recurrent|recurrent breast cancer_C0438105
C0438105|T047|ca br recurrence|recurrent breast cancer_C0438105
C0438105|T047|ca br recur|recurrent breast cancer_C0438105
C0438105|T047|ca br progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent brca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast ca|recurrent breast cancer_C0438105
C0438105|T047|breastca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breastca reoccur|recurrent breast cancer_C0438105
C0438105|T047|breastca recurrent|recurrent breast cancer_C0438105
C0438105|T047|breastca recurrence|recurrent breast cancer_C0438105
C0438105|T047|breastca recur|recurrent breast cancer_C0438105
C0438105|T047|breastca progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent breast adenocarc|recurrent breast cancer_C0438105
C0438105|T047|breastca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|ca ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|br cancer recurrence|recurrent breast cancer_C0438105
C0438105|T047|br cancer recur|recurrent breast cancer_C0438105
C0438105|T047|br cancer progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br cancer recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|br ca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br ca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br ca reoccur|recurrent breast cancer_C0438105
C0438105|T047|br ca recurrent|recurrent breast cancer_C0438105
C0438105|T047|br ca recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast recur|recurrent breast cancer_C0438105
C0438105|T047|br ca recur|recurrent breast cancer_C0438105
C0438105|T047|br cancer reoccur|recurrent breast cancer_C0438105
C0438105|T047|br cancer reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|br carc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br cancer reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br carc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br carc recurrent|recurrent breast cancer_C0438105
C0438105|T047|br carc recurrence|recurrent breast cancer_C0438105
C0438105|T047|br carc recur|recurrent breast cancer_C0438105
C0438105|T047|br carc progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma br recurrence|recurrent breast cancer_C0438105
C0438105|T047|br carc reoccur|recurrent breast cancer_C0438105
C0438105|T047|br carcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br ca progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc reoccur|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc recurrent|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc recurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc recur|recurrent breast cancer_C0438105
C0438105|T047|br adenocarc progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenoca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br adenoca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenoca reoccur|recurrent breast cancer_C0438105
C0438105|T047|br adenoca recurrent|recurrent breast cancer_C0438105
C0438105|T047|br adenoca recurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenoca recur|recurrent breast cancer_C0438105
C0438105|T047|br adenoca progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma recurrent|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma recur|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarcinoma ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|br adenocarcinoma reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma recurrence|recurrent breast cancer_C0438105
C0438105|T047|br malig progressive|recurrent breast cancer_C0438105
C0438105|T047|br malig recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca recur|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca progressive|recurrent breast cancer_C0438105
C0438105|T047|brca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|brca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|brca reoccur|recurrent breast cancer_C0438105
C0438105|T047|brca recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca recurrent|recurrent breast cancer_C0438105
C0438105|T047|brca recurrence|recurrent breast cancer_C0438105
C0438105|T047|brca progressive|recurrent breast cancer_C0438105
C0438105|T047|br tumor reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br tumor reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br tumor reoccur|recurrent breast cancer_C0438105
C0438105|T047|br tumor recurrent|recurrent breast cancer_C0438105
C0438105|T047|br tumor recurrence|recurrent breast cancer_C0438105
C0438105|T047|br tumor recur|recurrent breast cancer_C0438105
C0438105|T047|brca recur|recurrent breast cancer_C0438105
C0438105|T047|br tumor progressive|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarcinoma progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal recur|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast adenoca reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc reoccur|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc recurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc recurrence|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc recur|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc progressive|recurrent breast cancer_C0438105
C0438105|T047|adenocarc ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|breast adenocarc reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br malig recur|recurrent breast cancer_C0438105
C0438105|T047|tumor br progressive|recurrent breast cancer_C0438105
C0438105|T047|tumor br recurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br malignancy reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br malignancy reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal recur|recurrent breast cancer_C0438105
C0438105|T047|br malignancy reoccur|recurrent breast cancer_C0438105
C0438105|T047|br malignancy recurrence|recurrent breast cancer_C0438105
C0438105|T047|br malignancy recur|recurrent breast cancer_C0438105
C0438105|T047|br malignancy progressive|recurrent breast cancer_C0438105
C0438105|T047|br malig reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|br malig reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|br malig reoccur|recurrent breast cancer_C0438105
C0438105|T047|br malig recurrent|recurrent breast cancer_C0438105
C0438105|T047|br malignancy recurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor br recur|recurrent breast cancer_C0438105
C0438105|T047|tumor ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor br recurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor br reoccur|recurrent breast cancer_C0438105
C0438105|T047|tumor br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor breast progressive|recurrent breast cancer_C0438105
C0438105|T047|tumor breast recur|recurrent breast cancer_C0438105
C0438105|T047|tumor breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl recur|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|tumor dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|tumor breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|ca ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|ca ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br ca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast malig|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br cancer|recurrent breast cancer_C0438105
C0438105|T047|ca ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br malig|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence brca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence br carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breastca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal carc|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal malig|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|adenoca br progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl malig|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl carcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl carc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl cancer|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl ca|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence dctl adenocarc|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal cancer|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|cancer breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|cancer breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer breast recur|recurrent breast cancer_C0438105
C0438105|T047|adenoca br reoccur|recurrent breast cancer_C0438105
C0438105|T047|cancer br progressive|recurrent breast cancer_C0438105
C0438105|T047|cancer breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer br recur|recurrent breast cancer_C0438105
C0438105|T047|cancer br recurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer br reoccur|recurrent breast cancer_C0438105
C0438105|T047|cancer br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|adenoca br recurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer breast progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca br recurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer br recurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl recur|recurrent breast cancer_C0438105
C0438105|T047|adenoca br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal recur|recurrent breast cancer_C0438105
C0438105|T047|cancer ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast adenocarc|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast ca|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast recur|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast progressive|recurrent breast cancer_C0438105
C0438105|T047|adenoca br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|cancer dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence breast cancer|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal ca|recurrent breast cancer_C0438105
C0438105|T047|adenoca br recur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal ca|recurrent breast cancer_C0438105
C0438105|T047|carc dctl reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carc br progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast tumor|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal tumor|recurrent breast cancer_C0438105
C0438105|T047|carc dctl reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccur breastca|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal carcinoma|recurrent breast cancer_C0438105
C0438105|T047|carc ductal progressive|recurrent breast cancer_C0438105
C0438105|T047|carc ductal recur|recurrent breast cancer_C0438105
C0438105|T047|carc br reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl cancer|recurrent breast cancer_C0438105
C0438105|T047|carc ductal recurrence|recurrent breast cancer_C0438105
C0438105|T047|carc dctl reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl carc|recurrent breast cancer_C0438105
C0438105|T047|carc dctl recurrent|recurrent breast cancer_C0438105
C0438105|T047|carc dctl recur|recurrent breast cancer_C0438105
C0438105|T047|carc br recurrent|recurrent breast cancer_C0438105
C0438105|T047|carc br recurrence|recurrent breast cancer_C0438105
C0438105|T047|carc br reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|carc breast progressive|recurrent breast cancer_C0438105
C0438105|T047|carc breast recur|recurrent breast cancer_C0438105
C0438105|T047|carc breast recurrence|recurrent breast cancer_C0438105
C0438105|T047|carc breast recurrent|recurrent breast cancer_C0438105
C0438105|T047|carc breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|carc breast reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carc br recur|recurrent breast cancer_C0438105
C0438105|T047|carc breast reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|carc dctl progressive|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal malig|recurrent breast cancer_C0438105
C0438105|T047|carc dctl recurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal carc|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl ca|recurrent breast cancer_C0438105
C0438105|T047|carc ductal reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br adenoca|recurrent breast cancer_C0438105
C0438105|T047|carc ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccur breast malig|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccurrent br adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl carcinoma|recurrent breast cancer_C0438105
C0438105|T047|adenoca breast reoccur|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl malignancy|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl tumor|recurrent breast cancer_C0438105
C0438105|T047|ca ductal reoccurrent|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal adenoca|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal adenocarc|recurrent breast cancer_C0438105
C0438105|T047|reoccur ductal adenocarcinoma|recurrent breast cancer_C0438105
C0438105|T047|reoccur dctl malig|recurrent breast cancer_C0438105
C0438105|T047|carc ductal recurrent|recurrent breast cancer_C0438105
C0438105|T047|carc br reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|carc ductal reoccurrence|recurrent breast cancer_C0438105
C0438105|T047|reoccurrence ductal cancer|recurrent breast cancer_C0438105
C0438106|T047|recurrent metastasis|metastatic recurrence_C0438106
C0438106|T047|reoccurrent spread|metastatic recurrence_C0438106
C0438106|T047|distant recurrence|metastatic recurrence_C0438106
C0438106|T047|reoccurrent metastatic|metastatic recurrence_C0438106
C0438106|T047|reoccurrent metastasize|metastatic recurrence_C0438106
C0438106|T047|reoccurrent metastasis|metastatic recurrence_C0438106
C0438106|T047|reoccurrent metastases|metastatic recurrence_C0438106
C0438106|T047|metastatic recur|metastatic recurrence_C0438106
C0438106|T047|metastatic progressive|metastatic recurrence_C0438106
C0438106|T047|reoccurrent met|metastatic recurrence_C0438106
C0438106|T047|reoccurrent mediastatic|metastatic recurrence_C0438106
C0438106|T047|disseminated progressive|metastatic recurrence_C0438106
C0438106|T047|disseminated reoccurrent|metastatic recurrence_C0438106
C0438106|T047|disseminated reoccurrence|metastatic recurrence_C0438106
C0438106|T047|disseminated reoccur|metastatic recurrence_C0438106
C0438106|T047|recurrent spread|metastatic recurrence_C0438106
C0438106|T047|recurrent disseminated|metastatic recurrence_C0438106
C0438106|T047|recurrent metastatic|metastatic recurrence_C0438106
C0438106|T047|disseminated recurrent|metastatic recurrence_C0438106
C0438106|T047|disseminated recurrence|metastatic recurrence_C0438106
C0438106|T047|recurrent mediastatic|metastatic recurrence_C0438106
C0438106|T047|recurrent met|metastatic recurrence_C0438106
C0438106|T047|recurrent metastases|metastatic recurrence_C0438106
C0438106|T047|recurrent metastasize|metastatic recurrence_C0438106
C0438106|T047|disseminated recur|metastatic recurrence_C0438106
C0438106|T047|met recur|metastatic recurrence_C0438106
C0438106|T047|mediastatic recur|metastatic recurrence_C0438106
C0438106|T047|metastasize recurrence|metastatic recurrence_C0438106
C0438106|T047|metastasize recur|metastatic recurrence_C0438106
C0438106|T047|metastasize progressive|metastatic recurrence_C0438106
C0438106|T047|metastasis reoccurrent|metastatic recurrence_C0438106
C0438106|T047|metastasis reoccur|metastatic recurrence_C0438106
C0438106|T047|metastasis recurrent|metastatic recurrence_C0438106
C0438106|T047|metastasis recurrence|metastatic recurrence_C0438106
C0438106|T047|metastasis recur|metastatic recurrence_C0438106
C0438106|T047|metastasis progressive|metastatic recurrence_C0438106
C0438106|T047|spread progressive|metastatic recurrence_C0438106
C0438106|T047|spread recur|metastatic recurrence_C0438106
C0438106|T047|metastasize recurrent|metastatic recurrence_C0438106
C0438106|T047|metastases reoccurrent|metastatic recurrence_C0438106
C0438106|T047|metastases reoccur|metastatic recurrence_C0438106
C0438106|T047|metastases recurrent|metastatic recurrence_C0438106
C0438106|T047|metastases recurrence|metastatic recurrence_C0438106
C0438106|T047|metastases recur|metastatic recurrence_C0438106
C0438106|T047|spread recurrence|metastatic recurrence_C0438106
C0438106|T047|spread recurrent|metastatic recurrence_C0438106
C0438106|T047|spread reoccur|metastatic recurrence_C0438106
C0438106|T047|spread reoccurrence|metastatic recurrence_C0438106
C0438106|T047|metastases progressive|metastatic recurrence_C0438106
C0438106|T047|spread reoccurrent|metastatic recurrence_C0438106
C0438106|T047|reoccur disseminated|metastatic recurrence_C0438106
C0438106|T047|metastases reoccurrence|metastatic recurrence_C0438106
C0438106|T047|metastasize reoccur|metastatic recurrence_C0438106
C0438106|T047|metastasize reoccurrence|metastatic recurrence_C0438106
C0438106|T047|metastasize reoccurrent|metastatic recurrence_C0438106
C0438106|T047|mediastatic recurrence|metastatic recurrence_C0438106
C0438106|T047|mediastatic recurrent|metastatic recurrence_C0438106
C0438106|T047|mediastatic reoccur|metastatic recurrence_C0438106
C0438106|T047|mediastatic reoccurrence|metastatic recurrence_C0438106
C0438106|T047|mediastatic reoccurrent|metastatic recurrence_C0438106
C0438106|T047|met progressive|metastatic recurrence_C0438106
C0438106|T047|met recurrence|metastatic recurrence_C0438106
C0438106|T047|met recurrent|metastatic recurrence_C0438106
C0438106|T047|met reoccurrence|metastatic recurrence_C0438106
C0438106|T047|reoccur spread|metastatic recurrence_C0438106
C0438106|T047|recurrence disseminated|metastatic recurrence_C0438106
C0438106|T047|reoccur metastatic|metastatic recurrence_C0438106
C0438106|T047|reoccur metastasize|metastatic recurrence_C0438106
C0438106|T047|met reoccurrent|metastatic recurrence_C0438106
C0438106|T047|reoccur metastasis|metastatic recurrence_C0438106
C0438106|T047|recurrence mediastatic|metastatic recurrence_C0438106
C0438106|T047|recurrence met|metastatic recurrence_C0438106
C0438106|T047|recurrence metastases|metastatic recurrence_C0438106
C0438106|T047|recurrence metastasis|metastatic recurrence_C0438106
C0438106|T047|recurrence metastasize|metastatic recurrence_C0438106
C0438106|T047|recurrence metastatic|metastatic recurrence_C0438106
C0438106|T047|recurrence spread|metastatic recurrence_C0438106
C0438106|T047|reoccur metastases|metastatic recurrence_C0438106
C0438106|T047|reoccur met|metastatic recurrence_C0438106
C0438106|T047|reoccur mediastatic|metastatic recurrence_C0438106
C0438106|T047|mediastatic progressive|metastatic recurrence_C0438106
C0438106|T047|metastasis reoccurrence|metastatic recurrence_C0438106
C0438106|T047|met reoccur|metastatic recurrence_C0438106
C0438106|T047|recur metastases|metastatic recurrence_C0438106
C0438106|T047|metastatic reoccurrence|metastatic recurrence_C0438106
C0438106|T047|metastatic reoccurrent|metastatic recurrence_C0438106
C0438106|T047|reoccurrent disseminated|metastatic recurrence_C0438106
C0438106|T047|progressive metastasize|metastatic recurrence_C0438106
C0438106|T047|reoccurrence spread|metastatic recurrence_C0438106
C0438106|T047|reoccurrence metastatic|metastatic recurrence_C0438106
C0438106|T047|reoccurrence metastasize|metastatic recurrence_C0438106
C0438106|T047|reoccurrence metastasis|metastatic recurrence_C0438106
C0438106|T047|reoccurrence metastases|metastatic recurrence_C0438106
C0438106|T047|recur mediastatic|metastatic recurrence_C0438106
C0438106|T047|reoccurrence met|metastatic recurrence_C0438106
C0438106|T047|reoccurrence mediastatic|metastatic recurrence_C0438106
C0438106|T047|progressive mediastatic|metastatic recurrence_C0438106
C0438106|T047|progressive metastatic|metastatic recurrence_C0438106
C0438106|T047|progressive spread|metastatic recurrence_C0438106
C0438106|T047|recur metastatic|metastatic recurrence_C0438106
C0438106|T047|metastatic reoccur|metastatic recurrence_C0438106
C0438106|T047|recur met|metastatic recurrence_C0438106
C0438106|T047|progressive metastases|metastatic recurrence_C0438106
C0438106|T047|recur spread|metastatic recurrence_C0438106
C0438106|T047|progressive disseminated|metastatic recurrence_C0438106
C0438106|T047|progressive metastasis|metastatic recurrence_C0438106
C0438106|T047|reoccurrence disseminated|metastatic recurrence_C0438106
C0438106|T047|recur metastasis|metastatic recurrence_C0438106
C0438106|T047|recur disseminated|metastatic recurrence_C0438106
C0438106|T047|progressive met|metastatic recurrence_C0438106
C0438106|T047|metastatic recurrence|metastatic recurrence_C0438106
C0438106|T047|recur metastasize|metastatic recurrence_C0438106
C0438106|T047|metastatic recurrent|metastatic recurrence_C0438106
C0438110|T047|ductal reoccurrence|recurrent breast_C0438110
C0438110|T047|br recurrence|recurrent breast_C0438110
C0438110|T047|breast reoccurrent|recurrent breast_C0438110
C0438110|T047|recur breast|recurrent breast_C0438110
C0438110|T047|recurrence dctl|recurrent breast_C0438110
C0438110|T047|in-breast recurrence|recurrent breast_C0438110
C0438110|T047|dctl recurrence|recurrent breast_C0438110
C0438110|T047|reoccurrent dctl|recurrent breast_C0438110
C0438110|T047|progressive breast|recurrent breast_C0438110
C0438110|T047|dctl reoccurrent|recurrent breast_C0438110
C0438110|T047|recurrent ductal|recurrent breast_C0438110
C0438110|T047|reoccurrent breast|recurrent breast_C0438110
C0438110|T047|ductal recurrence|recurrent breast_C0438110
C0438110|T047|br recur|recurrent breast_C0438110
C0438110|T047|dctl reoccurrence|recurrent breast_C0438110
C0438110|T047|recurrence breast|recurrent breast_C0438110
C0438110|T047|reoccurrence br|recurrent breast_C0438110
C0438110|T047|dctl recur|recurrent breast_C0438110
C0438110|T047|dctl reoccur|recurrent breast_C0438110
C0438110|T047|ductal recurrent|recurrent breast_C0438110
C0438110|T047|recur ductal|recurrent breast_C0438110
C0438110|T047|recurrent dctl|recurrent breast_C0438110
C0438110|T047|recurrence br|recurrent breast_C0438110
C0438110|T047|recur br|recurrent breast_C0438110
C0438110|T047|ductal progressive|recurrent breast_C0438110
C0438110|T047|br progressive|recurrent breast_C0438110
C0438110|T047|reoccurrence breast|recurrent breast_C0438110
C0438110|T047|progressive dctl|recurrent breast_C0438110
C0438110|T047|recurrence ductal|recurrent breast_C0438110
C0438110|T047|ductal reoccur|recurrent breast_C0438110
C0438110|T047|dctl recurrent|recurrent breast_C0438110
C0438110|T047|reoccur ductal|recurrent breast_C0438110
C0438110|T047|recurrent br|recurrent breast_C0438110
C0438110|T047|reoccur dctl|recurrent breast_C0438110
C0438110|T047|dctl progressive|recurrent breast_C0438110
C0438110|T047|reoccur breast|recurrent breast_C0438110
C0438110|T047|progressive ductal|recurrent breast_C0438110
C0438110|T047|reoccurrence dctl|recurrent breast_C0438110
C0438110|T047|recur dctl|recurrent breast_C0438110
C0438110|T047|breast recurrence|recurrent breast_C0438110
C0438110|T047|br reoccurrent|recurrent breast_C0438110
C0438110|T047|recurrent breast|recurrent breast_C0438110
C0438110|T047|breast recurrent|recurrent breast_C0438110
C0438110|T047|breast reoccur|recurrent breast_C0438110
C0438110|T047|reoccurrent ductal|recurrent breast_C0438110
C0438110|T047|reoccurrence ductal|recurrent breast_C0438110
C0438110|T047|breast reoccurrence|recurrent breast_C0438110
C0438110|T047|br reoccurrence|recurrent breast_C0438110
C0438110|T047|breast recur|recurrent breast_C0438110
C0438110|T047|progressive br|recurrent breast_C0438110
C0438110|T047|br reoccur|recurrent breast_C0438110
C0438110|T047|reoccurrent br|recurrent breast_C0438110
C0438110|T047|br recurrent|recurrent breast_C0438110
C0438110|T047|reoccur br|recurrent breast_C0438110
C0438110|T047|ductal recur|recurrent breast_C0438110
C0438110|T047|breast progressive|recurrent breast_C0438110
C0438110|T047|ductal reoccurrent|recurrent breast_C0438110
C0438111|T047|recurrent breast spread|recurrent breast metastatic_C0438111
C0438111|T047|recur breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast recur|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|recur breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recur breast spread|recurrent breast metastatic_C0438111
C0438111|T047|recur breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recur breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|metastases br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastases br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|metastases br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastases br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastases br progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastases br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastases br recur|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastases breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recur breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br met|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|recur br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recur breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|metastases dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|recur br spread|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recur br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recur br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastases ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|reoccur dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|recur br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recur br met|recurrent breast metastatic_C0438111
C0438111|T047|recur br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recur breast met|recurrent breast metastatic_C0438111
C0438111|T047|recur br metastases|recurrent breast metastatic_C0438111
C0438111|T047|met br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|met ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal met|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal met|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl met|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br progressive|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br recur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccur br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast recur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|met ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrent dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|met br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|met br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|met br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|met br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|met breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|met breast recur|recurrent breast metastatic_C0438111
C0438111|T047|met breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|met breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|met breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|met breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|met br recur|recurrent breast metastatic_C0438111
C0438111|T047|met breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|met dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|met dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|met dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|met dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|met dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|met dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|met ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|met ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|met ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|met ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|met ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|met dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|met br progressive|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl met|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccur breast spread|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal met|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recur ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recur dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|mediastatic dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast recur|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast met|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br met|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence br spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|spread breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|recurrence dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast metastasis|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast metastases|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast recur|recurrent breast metastatic_C0438111
C0438111|T047|recurrence breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|progressive breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|spread breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal met|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl met|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread breast recur|recurrent breast metastatic_C0438111
C0438111|T047|spread breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|progressive br spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|spread br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|spread br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br metastases|recurrent breast metastatic_C0438111
C0438111|T047|progressive br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|progressive br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|progressive br metastases|recurrent breast metastatic_C0438111
C0438111|T047|progressive br met|recurrent breast metastatic_C0438111
C0438111|T047|progressive br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|spread br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread br recur|recurrent breast metastatic_C0438111
C0438111|T047|spread br progressive|recurrent breast metastatic_C0438111
C0438111|T047|progressive br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastatic breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|recurrence br met|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br metastases|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal metastases|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccur ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrent breast disseminated|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasis dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasis ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br disseminated|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl metastatic|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl metastasize|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|spread dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence breast spread|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl metastasis|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl metastases|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl met|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal spread|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal metastatic|recurrent breast metastatic_C0438111
C0438111|T047|progressive dctl mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal metastasis|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br recur|recurrent breast metastatic_C0438111
C0438111|T047|metastatic br progressive|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br met|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br metastases|recurrent breast metastatic_C0438111
C0438111|T047|metastasize dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|metastasize ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal met|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal met|recurrent breast metastatic_C0438111
C0438111|T047|progressive ductal disseminated|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br spread|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrence dctl disseminated|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br spread|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|spread ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br metastasize|recurrent breast metastatic_C0438111
C0438111|T047|recurrent br metastasis|recurrent breast metastatic_C0438111
C0438111|T047|reoccurrent br metastatic|recurrent breast metastatic_C0438111
C0438111|T047|recurrence ductal metastasize|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive metastasize|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|br recur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br recur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br recur metastases|recurrent breast metastatic_C0438111
C0438111|T047|br recur met|recurrent breast metastatic_C0438111
C0438111|T047|br recur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br recur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br recur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br progressive spread|recurrent breast metastatic_C0438111
C0438111|T047|br progressive metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br progressive metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br progressive metastases|recurrent breast metastatic_C0438111
C0438111|T047|br progressive met|recurrent breast metastatic_C0438111
C0438111|T047|br progressive mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br progressive disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br progressive metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br recur spread|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent met|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br recurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|br recurrence met|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur met|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br progressive|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive metastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive met|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br recur|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br recurrence|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br recurrent|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence met|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent met|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent met|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br reoccur|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur met|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent met|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive met|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur met|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence met|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive disseminated|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast progressive mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence met|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur metastases|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur spread|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent met|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence met|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur spread|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|br reoccur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur metastases|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|br reoccurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur met|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|dctl recurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl reoccurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|dctl recur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|disseminated br reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur spread|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur met|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal recur|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast recur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent met|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence met|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast recur spread|recurrent breast metastatic_C0438111
C0438111|T047|breast recur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast recur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence met|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal progressive|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl reoccur|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur metastasize|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl recurrent|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl recurrence|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl recur|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur spread|recurrent breast metastatic_C0438111
C0438111|T047|disseminated dctl progressive|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence met|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur met|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|ductal recur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent met|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|breast reoccurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|breast recur metastasis|recurrent breast metastatic_C0438111
C0438111|T047|breast recurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|breast recur met|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent metastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive metastasis|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent metastasize|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent metastasis|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast recur|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast progressive|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence metastases|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent met|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence metastasis|recurrent breast metastatic_C0438111
C0438111|T047|dctl progressive disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence metastasize|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrent spread|recurrent breast metastatic_C0438111
C0438111|T047|ductal recurrence metastatic|recurrent breast metastatic_C0438111
C0438111|T047|breast recur mediastatic|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal reoccurrent|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|breast recur metastases|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal reoccur|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal recurrent|recurrent breast metastatic_C0438111
C0438111|T047|disseminated ductal recurrence|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive metastases|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast recurrence|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive met|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast reoccurrence|recurrent breast metastatic_C0438111
C0438111|T047|ductal reoccur disseminated|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive disseminated|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast recurrent|recurrent breast metastatic_C0438111
C0438111|T047|disseminated breast reoccur|recurrent breast metastatic_C0438111
C0438111|T047|ductal progressive mediastatic|recurrent breast metastatic_C0438111
C0438112|T047|reoccur adenoca|recurrent cancer_C0438112
C0438112|T047|progressive malignancy|recurrent cancer_C0438112
C0438112|T047|ca recur|recurrent cancer_C0438112
C0438112|T047|recurrent tumor|recurrent cancer_C0438112
C0438112|T047|reoccurrence malig|recurrent cancer_C0438112
C0438112|T047|progressive malig|recurrent cancer_C0438112
C0438112|T047|adenoca progressive|recurrent cancer_C0438112
C0438112|T047|adenocarc recurrent|recurrent cancer_C0438112
C0438112|T047|recurrent malig|recurrent cancer_C0438112
C0438112|T047|reoccurrence malignancy|recurrent cancer_C0438112
C0438112|T047|carc reoccurrent|recurrent cancer_C0438112
C0438112|T047|recur adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|cancer reoccur|recurrent cancer_C0438112
C0438112|T047|carcinoma reoccurrence|recurrent cancer_C0438112
C0438112|T047|reoccur adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|reoccur adenocarc|recurrent cancer_C0438112
C0438112|T047|recur adenocarc|recurrent cancer_C0438112
C0438112|T047|ca recurrent|recurrent cancer_C0438112
C0438112|T047|adenoca reoccurrent|recurrent cancer_C0438112
C0438112|T047|adenoca reoccurrence|recurrent cancer_C0438112
C0438112|T047|cancer reoccurrence|recurrent cancer_C0438112
C0438112|T047|ca recurrence|recurrent cancer_C0438112
C0438112|T047|carc reoccurrence|recurrent cancer_C0438112
C0438112|T047|ca recuring|recurrent cancer_C0438112
C0438112|T047|malig recur|recurrent cancer_C0438112
C0438112|T047|adenoca reoccur|recurrent cancer_C0438112
C0438112|T047|recurrent malignancy|recurrent cancer_C0438112
C0438112|T047|recur ca|recurrent cancer_C0438112
C0438112|T047|malig progressive|recurrent cancer_C0438112
C0438112|T047|reoccurrent ca|recurrent cancer_C0438112
C0438112|T047|progressive adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|ca progressive|recurrent cancer_C0438112
C0438112|T047|reoccurrence tumor|recurrent cancer_C0438112
C0438112|T047|reoccur cancer|recurrent cancer_C0438112
C0438112|T047|reoccur ca|recurrent cancer_C0438112
C0438112|T047|recurring cancer|recurrent cancer_C0438112
C0438112|T047|recurring ca|recurrent cancer_C0438112
C0438112|T047|recurring adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|recurring adenocarc|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recurrence|recurrent cancer_C0438112
C0438112|T047|recurring adenoca|recurrent cancer_C0438112
C0438112|T047|carc progressive|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recuring|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recur|recurrent cancer_C0438112
C0438112|T047|adenocarc recurring|recurrent cancer_C0438112
C0438112|T047|reoccurrent malig|recurrent cancer_C0438112
C0438112|T047|reoccurrent malignancy|recurrent cancer_C0438112
C0438112|T047|cancer reoccurrent|recurrent cancer_C0438112
C0438112|T047|progressive adenocarc|recurrent cancer_C0438112
C0438112|T047|progressive adenoca|recurrent cancer_C0438112
C0438112|T047|reoccurrent adenoca|recurrent cancer_C0438112
C0438112|T047|reoccurrent cancer|recurrent cancer_C0438112
C0438112|T047|reoccurrent carc|recurrent cancer_C0438112
C0438112|T047|recur carc|recurrent cancer_C0438112
C0438112|T047|recur carcinoma|recurrent cancer_C0438112
C0438112|T047|reoccurrent carcinoma|recurrent cancer_C0438112
C0438112|T047|progressive carcinoma|recurrent cancer_C0438112
C0438112|T047|progressive carc|recurrent cancer_C0438112
C0438112|T047|progressive cancer|recurrent cancer_C0438112
C0438112|T047|recur cancer|recurrent cancer_C0438112
C0438112|T047|reoccurrent tumor|recurrent cancer_C0438112
C0438112|T047|recur adenoca|recurrent cancer_C0438112
C0438112|T047|recurring carcinoma|recurrent cancer_C0438112
C0438112|T047|recurring carc|recurrent cancer_C0438112
C0438112|T047|reoccur carcinoma|recurrent cancer_C0438112
C0438112|T047|carc reoccur|recurrent cancer_C0438112
C0438112|T047|reoccur carc|recurrent cancer_C0438112
C0438112|T047|reoccurrent adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|reoccurrent adenocarc|recurrent cancer_C0438112
C0438112|T047|progressive ca|recurrent cancer_C0438112
C0438112|T047|malig recurrence|recurrent cancer_C0438112
C0438112|T047|progressive tumor|recurrent cancer_C0438112
C0438112|T047|malig reoccurrent|recurrent cancer_C0438112
C0438112|T047|malignancy recurrence|recurrent cancer_C0438112
C0438112|T047|adenocarc reoccurrence|recurrent cancer_C0438112
C0438112|T047|carcinoma recurrnet|recurrent cancer_C0438112
C0438112|T047|adenocarc recurrnet|recurrent cancer_C0438112
C0438112|T047|cancer recurring|recurrent cancer_C0438112
C0438112|T047|recurrence malignancy|recurrent cancer_C0438112
C0438112|T047|recurrence malig|recurrent cancer_C0438112
C0438112|T047|recuring cancer|recurrent cancer_C0438112
C0438112|T047|tumor recur|recurrent cancer_C0438112
C0438112|T047|tumor progressive|recurrent cancer_C0438112
C0438112|T047|carc recuring|recurrent cancer_C0438112
C0438112|T047|tumor recurrence|recurrent cancer_C0438112
C0438112|T047|malig reoccurrence|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recurrnet|recurrent cancer_C0438112
C0438112|T047|ca reoccurrent|recurrent cancer_C0438112
C0438112|T047|carc recur|recurrent cancer_C0438112
C0438112|T047|reoccurrence adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|reoccurrence adenocarc|recurrent cancer_C0438112
C0438112|T047|reoccurrence adenoca|recurrent cancer_C0438112
C0438112|T047|reoccur tumor|recurrent cancer_C0438112
C0438112|T047|recur tumor|recurrent cancer_C0438112
C0438112|T047|adenocarc reoccur|recurrent cancer_C0438112
C0438112|T047|cancer recurrence|recurrent cancer_C0438112
C0438112|T047|recuring carc|recurrent cancer_C0438112
C0438112|T047|cancer recurrent|recurrent cancer_C0438112
C0438112|T047|malignancy recurrent|recurrent cancer_C0438112
C0438112|T047|recuring ca|recurrent cancer_C0438112
C0438112|T047|recuring adenocarc|recurrent cancer_C0438112
C0438112|T047|reoccurrence ca|recurrent cancer_C0438112
C0438112|T047|adenoca recurrence|recurrent cancer_C0438112
C0438112|T047|reoccurrence cancer|recurrent cancer_C0438112
C0438112|T047|recuring adenoca|recurrent cancer_C0438112
C0438112|T047|reoccurrence carc|recurrent cancer_C0438112
C0438112|T047|reoccurrence carcinoma|recurrent cancer_C0438112
C0438112|T047|ca recurrnet|recurrent cancer_C0438112
C0438112|T047|ca reoccurrence|recurrent cancer_C0438112
C0438112|T047|carc recurrent|recurrent cancer_C0438112
C0438112|T047|cancer recurrnet|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma progressive|recurrent cancer_C0438112
C0438112|T047|malignancy recur|recurrent cancer_C0438112
C0438112|T047|tumor reoccurrent|recurrent cancer_C0438112
C0438112|T047|carc recurring|recurrent cancer_C0438112
C0438112|T047|adenoca recurrnet|recurrent cancer_C0438112
C0438112|T047|tumor reoccurrence|recurrent cancer_C0438112
C0438112|T047|cancer progressive|recurrent cancer_C0438112
C0438112|T047|carc recurrnet|recurrent cancer_C0438112
C0438112|T047|ca reoccur|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recurring|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma recurrent|recurrent cancer_C0438112
C0438112|T047|recur malignancy|recurrent cancer_C0438112
C0438112|T047|recur malig|recurrent cancer_C0438112
C0438112|T047|tumor reoccur|recurrent cancer_C0438112
C0438112|T047|tumor recurrent|recurrent cancer_C0438112
C0438112|T047|recurrnet adenoca|recurrent cancer_C0438112
C0438112|T047|recurrnet adenocarc|recurrent cancer_C0438112
C0438112|T047|malig reoccur|recurrent cancer_C0438112
C0438112|T047|recuring carcinoma|recurrent cancer_C0438112
C0438112|T047|carcinoma recurrence|recurrent cancer_C0438112
C0438112|T047|malignancy reoccurrence|recurrent cancer_C0438112
C0438112|T047|ca recurring|recurrent cancer_C0438112
C0438112|T047|carcinoma reoccurrent|recurrent cancer_C0438112
C0438112|T047|carcinoma recurrent|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma reoccur|recurrent cancer_C0438112
C0438112|T047|malignancy reoccur|recurrent cancer_C0438112
C0438112|T047|carcinoma reoccur|recurrent cancer_C0438112
C0438112|T047|carcinoma recurring|recurrent cancer_C0438112
C0438112|T047|adenocarc reoccurrent|recurrent cancer_C0438112
C0438112|T047|carc recurrence|recurrent cancer_C0438112
C0438112|T047|adenocarc recurrence|recurrent cancer_C0438112
C0438112|T047|recurrnet adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|adenocarc recuring|recurrent cancer_C0438112
C0438112|T047|adenoca recurring|recurrent cancer_C0438112
C0438112|T047|carcinoma progressive|recurrent cancer_C0438112
C0438112|T047|recurrent adenoca|recurrent cancer_C0438112
C0438112|T047|recurrent adenocarc|recurrent cancer_C0438112
C0438112|T047|recurrent adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|recurrent ca|recurrent cancer_C0438112
C0438112|T047|recurrent cancer|recurrent cancer_C0438112
C0438112|T047|malignancy progressive|recurrent cancer_C0438112
C0438112|T047|recurrent carc|recurrent cancer_C0438112
C0438112|T047|recurrent carcinoma|recurrent cancer_C0438112
C0438112|T047|recuring adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|adenoca recurrent|recurrent cancer_C0438112
C0438112|T047|adenocarc recur|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma reoccurrence|recurrent cancer_C0438112
C0438112|T047|adenocarc progressive|recurrent cancer_C0438112
C0438112|T047|recurrence carcinoma|recurrent cancer_C0438112
C0438112|T047|recurrence adenoca|recurrent cancer_C0438112
C0438112|T047|recurrence adenocarc|recurrent cancer_C0438112
C0438112|T047|recurrence adenocarcinoma|recurrent cancer_C0438112
C0438112|T047|adenocarcinoma reoccurrent|recurrent cancer_C0438112
C0438112|T047|carcinoma recur|recurrent cancer_C0438112
C0438112|T047|adenoca recuring|recurrent cancer_C0438112
C0438112|T047|cancer recuring|recurrent cancer_C0438112
C0438112|T047|recurrence ca|recurrent cancer_C0438112
C0438112|T047|recurrence cancer|recurrent cancer_C0438112
C0438112|T047|recurrence tumor|recurrent cancer_C0438112
C0438112|T047|reoccur malignancy|recurrent cancer_C0438112
C0438112|T047|recurrence carc|recurrent cancer_C0438112
C0438112|T047|recurrnet carcinoma|recurrent cancer_C0438112
C0438112|T047|reoccur malig|recurrent cancer_C0438112
C0438112|T047|adenoca recur|recurrent cancer_C0438112
C0438112|T047|malig recurrent|recurrent cancer_C0438112
C0438112|T047|cancer recur|recurrent cancer_C0438112
C0438112|T047|recurrnet carc|recurrent cancer_C0438112
C0438112|T047|carcinoma recuring|recurrent cancer_C0438112
C0438112|T047|recurrnet cancer|recurrent cancer_C0438112
C0438112|T047|malignancy reoccurrent|recurrent cancer_C0438112
C0438112|T047|recurrnet ca|recurrent cancer_C0438112
C0438113|T047|carc progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur met|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur met|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|recurrence met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|carc recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carc reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|recurrent mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|spread ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|tumor recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|tumor reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarc recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur met|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|ca progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur met|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccur spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|cancer recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|ca reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrence metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|spread adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|reoccurrent disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur met|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|adenoca recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|met tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|met malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur met|recurrent cancer metastatic_C0438113
C0438113|T047|malig recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastases adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasis carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy progressive spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recur spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malignancy reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|met carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|met carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|met cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|met ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur met|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|met carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|met malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|met carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|malig recurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|met malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccur spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|malig reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|met adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|mediastatic tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|met adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|adenocarcinoma recurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur met carc|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur met malig|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|recur met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recur met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recur met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur met ca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis malig|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasis tumor|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated tumor|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive disseminated adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive metastases adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met tumor|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met cancer|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|recur mediastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|progressive mediastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|progressive met ca|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic carc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur disseminated ca|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread malig|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenoca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize tumor progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread tumor|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent spread|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic tumor|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc progressive|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread adenoca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic malig|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread ca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread cancer|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread carc|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic carc|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic ca|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic adenocarcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarcinoma progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur spread carcinoma|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic adenocarc recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic cancer|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy recur|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic malignancy|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malignancy progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastatic adenocarc|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence spread|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence metastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence metastases|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence met|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence disseminated|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer progressive|recurrent cancer metastatic_C0438113
C0438113|T047|recur metastasize tumor|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic cancer reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize carcinoma recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrence mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastatic ca progressive|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent metastasize|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig reoccur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig recurrent|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig recurrence|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig recur|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig progressive|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent metastasis|recurrent cancer metastatic_C0438113
C0438113|T047|metastasize malig reoccurrence|recurrent cancer metastatic_C0438113
C0438113|T047|disseminated tumor reoccurrent|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent metastases|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent mediastatic|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent met|recurrent cancer metastatic_C0438113
C0438113|T047|carcinoma reoccurrent disseminated|recurrent cancer metastatic_C0438113
C0438120|T047|LF Breast Cancer Recurrence|recurrent breast cancer_C0438120
C0438120|T047|RT Breast Cancer Recurrence|recurrent breast cancer_C0438120
C0438204|T047|axillary recurrence|axillary recurrence_C0438204
C0441771|T047|stage III|stage IIIC_C0441771
C0441771|T047|stage 3|stage IIIC_C0441771
C0441771|T047|stage 3A|stage IIIC_C0441771
C0441771|T047|stage 3B|stage IIIC_C0441771
C0441771|T047|stage 3C|stage IIIC_C0441771
C0441771|T047|stage IIIB|stage IIIC_C0441771
C0441771|T047|stage IIIC|stage IIIC_C0441771
C0441771|T047|stage IIIA|stage IIIC_C0441771
C0441772|T047|stage IV|stage IV_C0441772
C0441772|T047|stage 4|stage IV_C0441772
C0441989|T047|Ipsilateral Recurrence|Ipsilateral Recurrence_C0441989
C0444498|T047|in-situ|intraductal_C0444498
C0444498|T047|intraductal|intraductal_C0444498
C0444498|T047|intraductl|intraductal_C0444498
C0444498|T047|in situ|intraductal_C0444498
C0500000|T047|positive axilla|positive lymph node_C0500000
C0500000|T047|metastatic axillary node|positive lymph node_C0500000
C0500000|T047|micrometastasis lymph node|positive lymph node_C0500000
C0500000|T047|positive lymph node|positive lymph node_C0500000
C0500000|T047|positive axillary node|positive lymph node_C0500000
C0500000|T047|metastatic lymph node|positive lymph node_C0500000
C0500000|T047|axillary nodal positive|positive lymph node_C0500000
C0500000|T047|axillary node metastatic|positive lymph node_C0500000
C0500000|T047|axillary node positive|positive lymph node_C0500000
C0500000|T047|lymph node metastatic|positive lymph node_C0500000
C0500000|T047|metastases to axilla|positive lymph node_C0500000
C0500000|T047|axillary nodal metastatic|positive lymph node_C0500000
C0500000|T047|metastases to axillary node|positive lymph node_C0500000
C0500000|T047|axillary nodal metastases|positive lymph node_C0500000
C0500000|T047|lymph node positive|positive lymph node_C0500000
C0500000|T047|metastases to lymph node|positive lymph node_C0500000
C0500000|T047|lymph node micrometastasis|positive lymph node_C0500000
C0684833|T192|CW Recurrence|CW Recurrence_C0684833
C0684833|T192|Recurrent Chest Wall Breast Cancer|CW Recurrence_C0684833
C0851238|T061|Lumpectomy|Lumpectomy_C0851238
C1134719|T047|infiltr breast ca|IDC_C1134719
C1134719|T047|infiltr breast adenocarcinoma|IDC_C1134719
C1134719|T047|infiltr breast adenocarc|IDC_C1134719
C1134719|T047|infiltr breast cancer|IDC_C1134719
C1134719|T047|infiltrduct lobular ca|IDC_C1134719
C1134719|T047|infiltr breast adenoca|IDC_C1134719
C1134719|T047|infil br carc|IDC_C1134719
C1134719|T047|infil br cancer|IDC_C1134719
C1134719|T047|infil br ca|IDC_C1134719
C1134719|T047|infil br adenocarcinoma|IDC_C1134719
C1134719|T047|infiltr breast carc|IDC_C1134719
C1134719|T047|infiltr br carcinoma|IDC_C1134719
C1134719|T047|infil lobular carc|IDC_C1134719
C1134719|T047|infiltr br cancer|IDC_C1134719
C1134719|T047|infiltr br ca|IDC_C1134719
C1134719|T047|infiltr br adenocarcinoma|IDC_C1134719
C1134719|T047|infiltr br adenocarc|IDC_C1134719
C1134719|T047|infiltr br adenoca|IDC_C1134719
C1134719|T047|infil lobular carcinoma|IDC_C1134719
C1134719|T047|infil lobular cancer|IDC_C1134719
C1134719|T047|infil lobular ca|IDC_C1134719
C1134719|T047|infil lobular adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating lobular carc|IDC_C1134719
C1134719|T047|infitrating lobular carcinoma|IDC_C1134719
C1134719|T047|infiltr br carc|IDC_C1134719
C1134719|T047|infil br adenocarc|IDC_C1134719
C1134719|T047|infiltrduct br adenocarc|IDC_C1134719
C1134719|T047|infiltrating lobular carc|IDC_C1134719
C1134719|T047|infiltrduct dctl ca|IDC_C1134719
C1134719|T047|infiltrduct lobular cancer|IDC_C1134719
C1134719|T047|infiltrduct dctl adenocarc|IDC_C1134719
C1134719|T047|infiltrduct dctl adenoca|IDC_C1134719
C1134719|T047|infiltrduct breast carcinoma|IDC_C1134719
C1134719|T047|infiltrduct breast carc|IDC_C1134719
C1134719|T047|infiltrduct breast cancer|IDC_C1134719
C1134719|T047|infiltrduct breast ca|IDC_C1134719
C1134719|T047|infiltrduct breast adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating ductal adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating ductal ca|IDC_C1134719
C1134719|T047|infitrating ductal cancer|IDC_C1134719
C1134719|T047|infitrating ductal carc|IDC_C1134719
C1134719|T047|infitrating ductal carcinoma|IDC_C1134719
C1134719|T047|infiltrduct breast adenocarc|IDC_C1134719
C1134719|T047|infiltrduct breast adenoca|IDC_C1134719
C1134719|T047|infiltrduct br carcinoma|IDC_C1134719
C1134719|T047|infiltrduct br carc|IDC_C1134719
C1134719|T047|infiltrduct br cancer|IDC_C1134719
C1134719|T047|infiltrduct br ca|IDC_C1134719
C1134719|T047|infiltrduct br adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating lobular adenoca|IDC_C1134719
C1134719|T047|infitrating lobular adenocarc|IDC_C1134719
C1134719|T047|infitrating lobular adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating lobular ca|IDC_C1134719
C1134719|T047|infitrating lobular cancer|IDC_C1134719
C1134719|T047|infil lobular adenocarc|IDC_C1134719
C1134719|T047|infiltrduct br adenoca|IDC_C1134719
C1134719|T047|infiltrating lobular carcinoma|IDC_C1134719
C1134719|T047|infil br adenoca|IDC_C1134719
C1134719|T047|infil lobular adenoca|IDC_C1134719
C1134719|T047|infil ductal adenocarcinoma|IDC_C1134719
C1134719|T047|infil ductal carc|IDC_C1134719
C1134719|T047|infltrtng breast ca|IDC_C1134719
C1134719|T047|infltrtng breast cancer|IDC_C1134719
C1134719|T047|infltrtng breast carc|IDC_C1134719
C1134719|T047|infltrtng breast carcinoma|IDC_C1134719
C1134719|T047|infltrtng dctl adenoca|IDC_C1134719
C1134719|T047|infltrtng dctl adenocarc|IDC_C1134719
C1134719|T047|infltrtng dctl adenocarcinoma|IDC_C1134719
C1134719|T047|infltrtng dctl ca|IDC_C1134719
C1134719|T047|infltrtng dctl cancer|IDC_C1134719
C1134719|T047|invasive br ca|IDC_C1134719
C1134719|T047|invasive br cancer|IDC_C1134719
C1134719|T047|invasive br carc|IDC_C1134719
C1134719|T047|infltrtng dctl carc|IDC_C1134719
C1134719|T047|infltrtng dctl carcinoma|IDC_C1134719
C1134719|T047|infltrtng ductal adenoca|IDC_C1134719
C1134719|T047|infltrtng ductal adenocarc|IDC_C1134719
C1134719|T047|infltrtng ductal adenocarcinoma|IDC_C1134719
C1134719|T047|infltrtng ductal ca|IDC_C1134719
C1134719|T047|infltrtng ductal cancer|IDC_C1134719
C1134719|T047|infltrtng ductal carc|IDC_C1134719
C1134719|T047|infltrtng ductal carcinoma|IDC_C1134719
C1134719|T047|infltrtng lobular adenoca|IDC_C1134719
C1134719|T047|infil dctl cancer|IDC_C1134719
C1134719|T047|infil dctl carc|IDC_C1134719
C1134719|T047|infil dctl carcinoma|IDC_C1134719
C1134719|T047|infil ductal adenoca|IDC_C1134719
C1134719|T047|infiltrating lobular ca|IDC_C1134719
C1134719|T047|infiltrating lobular adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrating lobular adenocarc|IDC_C1134719
C1134719|T047|infltrtng breast adenocarcinoma|IDC_C1134719
C1134719|T047|infltrtng breast adenocarc|IDC_C1134719
C1134719|T047|invasive br adenocarcinoma|IDC_C1134719
C1134719|T047|invasive br adenocarc|IDC_C1134719
C1134719|T047|infil ductal cancer|IDC_C1134719
C1134719|T047|infil ductal ca|IDC_C1134719
C1134719|T047|infiltrduct dctl cancer|IDC_C1134719
C1134719|T047|Multifocal IDC|IDC_C1134719
C1134719|T047|infiltrating lobular cancer|IDC_C1134719
C1134719|T047|infil ductal adenocarc|IDC_C1134719
C1134719|T047|infiltrating ductal carc|IDC_C1134719
C1134719|T047|infil br carcinoma|IDC_C1134719
C1134719|T047|infil breast adenoca|IDC_C1134719
C1134719|T047|infil breast adenocarc|IDC_C1134719
C1134719|T047|infil breast adenocarcinoma|IDC_C1134719
C1134719|T047|infil breast ca|IDC_C1134719
C1134719|T047|infil breast cancer|IDC_C1134719
C1134719|T047|infil breast carc|IDC_C1134719
C1134719|T047|infil ductal carcinoma|IDC_C1134719
C1134719|T047|infiltrating ductal carcinoma|IDC_C1134719
C1134719|T047|infil dctl adenoca|IDC_C1134719
C1134719|T047|infil dctl adenocarc|IDC_C1134719
C1134719|T047|infltrtng br adenoca|IDC_C1134719
C1134719|T047|infltrtng br adenocarc|IDC_C1134719
C1134719|T047|infltrtng br adenocarcinoma|IDC_C1134719
C1134719|T047|infltrtng br ca|IDC_C1134719
C1134719|T047|infltrtng br cancer|IDC_C1134719
C1134719|T047|infltrtng br carc|IDC_C1134719
C1134719|T047|infltrtng br carcinoma|IDC_C1134719
C1134719|T047|infltrtng breast adenoca|IDC_C1134719
C1134719|T047|infil dctl adenocarcinoma|IDC_C1134719
C1134719|T047|infil dctl ca|IDC_C1134719
C1134719|T047|infiltrating lobular adenoca|IDC_C1134719
C1134719|T047|invasive br adenoca|IDC_C1134719
C1134719|T047|infil breast carcinoma|IDC_C1134719
C1134719|T047|infiltrating ductal cancer|IDC_C1134719
C1134719|T047|infiltrduct dctl adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating ductal adenoca|IDC_C1134719
C1134719|T047|invasive ductal cancer|IDC_C1134719
C1134719|T047|invasive ductal ca|IDC_C1134719
C1134719|T047|infitrating breast ca|IDC_C1134719
C1134719|T047|invasive ductal adenocarcinoma|IDC_C1134719
C1134719|T047|invasive ductal adenocarc|IDC_C1134719
C1134719|T047|infiltrduct ductal adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrduct ductal adenocarc|IDC_C1134719
C1134719|T047|infiltrduct ductal adenoca|IDC_C1134719
C1134719|T047|infitrating breast cancer|IDC_C1134719
C1134719|T047|infitrating breast carc|IDC_C1134719
C1134719|T047|infiltrduct dctl carcinoma|IDC_C1134719
C1134719|T047|infiltrduct dctl carc|IDC_C1134719
C1134719|T047|invasive dctl adenoca|IDC_C1134719
C1134719|T047|invasive ductal carc|IDC_C1134719
C1134719|T047|invasive breast carcinoma|IDC_C1134719
C1134719|T047|infiltrating br carcinoma|IDC_C1134719
C1134719|T047|infiltrating breast adenoca|IDC_C1134719
C1134719|T047|infiltrating breast adenocarc|IDC_C1134719
C1134719|T047|infiltrating breast adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrating breast ca|IDC_C1134719
C1134719|T047|infiltrating breast cancer|IDC_C1134719
C1134719|T047|infiltrating breast carc|IDC_C1134719
C1134719|T047|infiltrating br adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating ductal adenocarc|IDC_C1134719
C1134719|T047|infiltrating br adenocarc|IDC_C1134719
C1134719|T047|infiltrating br adenoca|IDC_C1134719
C1134719|T047|infiltr lobular carcinoma|IDC_C1134719
C1134719|T047|infiltr lobular carc|IDC_C1134719
C1134719|T047|infiltrating br carc|IDC_C1134719
C1134719|T047|infiltrduct ductal ca|IDC_C1134719
C1134719|T047|invasive ductal carcinoma|IDC_C1134719
C1134719|T047|infiltrduct ductal cancer|IDC_C1134719
C1134719|T047|invasive dctl adenocarc|IDC_C1134719
C1134719|T047|invasive dctl adenocarcinoma|IDC_C1134719
C1134719|T047|invasive dctl ca|IDC_C1134719
C1134719|T047|infiltrduct lobular carc|IDC_C1134719
C1134719|T047|infiltrduct lobular carcinoma|IDC_C1134719
C1134719|T047|infitrating br adenoca|IDC_C1134719
C1134719|T047|infitrating br adenocarc|IDC_C1134719
C1134719|T047|infitrating br adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating br ca|IDC_C1134719
C1134719|T047|infitrating br cancer|IDC_C1134719
C1134719|T047|infitrating br carc|IDC_C1134719
C1134719|T047|infitrating br carcinoma|IDC_C1134719
C1134719|T047|infitrating breast adenoca|IDC_C1134719
C1134719|T047|infitrating breast adenocarc|IDC_C1134719
C1134719|T047|infitrating breast adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrating br cancer|IDC_C1134719
C1134719|T047|infiltrating br ca|IDC_C1134719
C1134719|T047|infiltrduct lobular adenocarcinoma|IDC_C1134719
C1134719|T047|invasive lobular carcinoma|IDC_C1134719
C1134719|T047|invasive lobular carc|IDC_C1134719
C1134719|T047|invasive lobular cancer|IDC_C1134719
C1134719|T047|invasive lobular ca|IDC_C1134719
C1134719|T047|invasive lobular adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrduct lobular adenocarc|IDC_C1134719
C1134719|T047|infiltrduct lobular adenoca|IDC_C1134719
C1134719|T047|invasive lobular adenocarc|IDC_C1134719
C1134719|T047|invasive lobular adenoca|IDC_C1134719
C1134719|T047|infiltrduct ductal carcinoma|IDC_C1134719
C1134719|T047|infiltrduct ductal carc|IDC_C1134719
C1134719|T047|infiltr lobular cancer|IDC_C1134719
C1134719|T047|infiltr lobular ca|IDC_C1134719
C1134719|T047|infiltr ductal carcinoma|IDC_C1134719
C1134719|T047|infiltrating breast carcinoma|IDC_C1134719
C1134719|T047|infiltrating dctl carcinoma|IDC_C1134719
C1134719|T047|infiltrating dctl carc|IDC_C1134719
C1134719|T047|infiltr ductal adenoca|IDC_C1134719
C1134719|T047|infiltr dctl carcinoma|IDC_C1134719
C1134719|T047|infiltr dctl carc|IDC_C1134719
C1134719|T047|infiltrating dctl cancer|IDC_C1134719
C1134719|T047|infiltr dctl cancer|IDC_C1134719
C1134719|T047|infiltrating dctl ca|IDC_C1134719
C1134719|T047|infiltr dctl ca|IDC_C1134719
C1134719|T047|infitrating dctl cancer|IDC_C1134719
C1134719|T047|invasive br carcinoma|IDC_C1134719
C1134719|T047|infiltrating ductal adenoca|IDC_C1134719
C1134719|T047|infiltr lobular adenocarcinoma|IDC_C1134719
C1134719|T047|invasive breast adenocarc|IDC_C1134719
C1134719|T047|infitrating dctl carc|IDC_C1134719
C1134719|T047|infitrating dctl carcinoma|IDC_C1134719
C1134719|T047|infiltr dctl adenocarcinoma|IDC_C1134719
C1134719|T047|infiltrating dctl adenoca|IDC_C1134719
C1134719|T047|infiltrating dctl adenocarc|IDC_C1134719
C1134719|T047|infltrtng lobular adenocarcinoma|IDC_C1134719
C1134719|T047|infltrtng lobular adenocarc|IDC_C1134719
C1134719|T047|infiltrating dctl adenocarcinoma|IDC_C1134719
C1134719|T047|invasive breast carc|IDC_C1134719
C1134719|T047|invasive breast cancer|IDC_C1134719
C1134719|T047|invasive breast adenoca|IDC_C1134719
C1134719|T047|invasive breast ca|IDC_C1134719
C1134719|T047|infiltr dctl adenocarc|IDC_C1134719
C1134719|T047|infiltr ductal adenocarc|IDC_C1134719
C1134719|T047|infiltr lobular adenocarc|IDC_C1134719
C1134719|T047|infiltr breast carcinoma|IDC_C1134719
C1134719|T047|infitrating breast carcinoma|IDC_C1134719
C1134719|T047|infiltr lobular adenoca|IDC_C1134719
C1134719|T047|infltrtng lobular carcinoma|IDC_C1134719
C1134719|T047|infltrtng lobular carc|IDC_C1134719
C1134719|T047|infltrtng lobular cancer|IDC_C1134719
C1134719|T047|infltrtng lobular ca|IDC_C1134719
C1134719|T047|infiltr ductal carc|IDC_C1134719
C1134719|T047|infiltrating ductal ca|IDC_C1134719
C1134719|T047|infiltr dctl adenoca|IDC_C1134719
C1134719|T047|infiltrating ductal adenocarcinoma|IDC_C1134719
C1134719|T047|invasive dctl carc|IDC_C1134719
C1134719|T047|invasive dctl carcinoma|IDC_C1134719
C1134719|T047|infiltr ductal cancer|IDC_C1134719
C1134719|T047|infiltr ductal ca|IDC_C1134719
C1134719|T047|invasive ductal adenoca|IDC_C1134719
C1134719|T047|infitrating dctl adenoca|IDC_C1134719
C1134719|T047|infitrating dctl adenocarc|IDC_C1134719
C1134719|T047|infitrating dctl adenocarcinoma|IDC_C1134719
C1134719|T047|infitrating dctl ca|IDC_C1134719
C1134719|T047|infiltrating ductal adenocarc|IDC_C1134719
C1134719|T047|infiltr ductal adenocarcinoma|IDC_C1134719
C1134719|T047|invasive dctl cancer|IDC_C1134719
C1134719|T047|invasive breast adenocarcinoma|IDC_C1134719
C1134720|T047|Recurrent IDC|Recurrent IDC_C1134720
C1268990|T047|breast|breast_C1268990
C1268990|T047|ductal|breast_C1268990
C1268990|T047|dctl|breast_C1268990
C1268990|T047|lobular|breast_C1268990
C1268990|T047|br|breast_C1268990
C1384494|T047|mediastatic carc|metastatic cancer_C1384494
C1384494|T047|mediastatic cancer|metastatic cancer_C1384494
C1384494|T047|mediastatic adenocarc|metastatic cancer_C1384494
C1384494|T047|malignancy metastatic|metastatic cancer_C1384494
C1384494|T047|malignancy metastasize|metastatic cancer_C1384494
C1384494|T047|malignancy metastasis|metastatic cancer_C1384494
C1384494|T047|malignancy metastases|metastatic cancer_C1384494
C1384494|T047|malignancy met|metastatic cancer_C1384494
C1384494|T047|adenocarc spread|metastatic cancer_C1384494
C1384494|T047|carcinoma spread|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma mediastatic|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma disseminated|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma met|metastatic cancer_C1384494
C1384494|T047|malignancy spread|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma spread|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma metastases|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma metastasize|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma metastatic|metastatic cancer_C1384494
C1384494|T047|mediastatic ca|metastatic cancer_C1384494
C1384494|T047|mediastatic adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|mediastatic adenoca|metastatic cancer_C1384494
C1384494|T047|adenocarcinoma metastasis|metastatic cancer_C1384494
C1384494|T047|metastasize carcinoma|metastatic cancer_C1384494
C1384494|T047|tumor spread|metastatic cancer_C1384494
C1384494|T047|adenoca metastasize|metastatic cancer_C1384494
C1384494|T047|adenoca metastatic|metastatic cancer_C1384494
C1384494|T047|metastasis adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|metastasis adenocarc|metastatic cancer_C1384494
C1384494|T047|metastasis adenoca|metastatic cancer_C1384494
C1384494|T047|metastases tumor|metastatic cancer_C1384494
C1384494|T047|metastases malignancy|metastatic cancer_C1384494
C1384494|T047|disseminated tumor|metastatic cancer_C1384494
C1384494|T047|cancer spread|metastatic cancer_C1384494
C1384494|T047|metastases malig|metastatic cancer_C1384494
C1384494|T047|malig disseminated|metastatic cancer_C1384494
C1384494|T047|malig mediastatic|metastatic cancer_C1384494
C1384494|T047|malig met|metastatic cancer_C1384494
C1384494|T047|malig metastases|metastatic cancer_C1384494
C1384494|T047|adenoca metastasis|metastatic cancer_C1384494
C1384494|T047|malig metastasis|metastatic cancer_C1384494
C1384494|T047|malig metastatic|metastatic cancer_C1384494
C1384494|T047|disseminated malignancy|metastatic cancer_C1384494
C1384494|T047|metastases carcinoma|metastatic cancer_C1384494
C1384494|T047|disseminated malig|metastatic cancer_C1384494
C1384494|T047|carc disseminated|metastatic cancer_C1384494
C1384494|T047|carc mediastatic|metastatic cancer_C1384494
C1384494|T047|carc met|metastatic cancer_C1384494
C1384494|T047|metastases carc|metastatic cancer_C1384494
C1384494|T047|carc metastases|metastatic cancer_C1384494
C1384494|T047|carc metastasis|metastatic cancer_C1384494
C1384494|T047|carc metastasize|metastatic cancer_C1384494
C1384494|T047|carc metastatic|metastatic cancer_C1384494
C1384494|T047|metastatic malig|metastatic cancer_C1384494
C1384494|T047|metastases cancer|metastatic cancer_C1384494
C1384494|T047|malig metastasize|metastatic cancer_C1384494
C1384494|T047|adenoca metastases|metastatic cancer_C1384494
C1384494|T047|adenoca met|metastatic cancer_C1384494
C1384494|T047|adenoca disseminated|metastatic cancer_C1384494
C1384494|T047|metastasize carc|metastatic cancer_C1384494
C1384494|T047|cancer metastatic|metastatic cancer_C1384494
C1384494|T047|cancer metastasize|metastatic cancer_C1384494
C1384494|T047|cancer metastasis|metastatic cancer_C1384494
C1384494|T047|cancer metastases|metastatic cancer_C1384494
C1384494|T047|cancer met|metastatic cancer_C1384494
C1384494|T047|cancer mediastatic|metastatic cancer_C1384494
C1384494|T047|cancer disseminated|metastatic cancer_C1384494
C1384494|T047|ca spread|metastatic cancer_C1384494
C1384494|T047|metastasize cancer|metastatic cancer_C1384494
C1384494|T047|metastasize ca|metastatic cancer_C1384494
C1384494|T047|metastasize adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|metastasize malig|metastatic cancer_C1384494
C1384494|T047|metastasize adenocarc|metastatic cancer_C1384494
C1384494|T047|metastasize malignancy|metastatic cancer_C1384494
C1384494|T047|metastasize adenoca|metastatic cancer_C1384494
C1384494|T047|metastasize tumor|metastatic cancer_C1384494
C1384494|T047|ca disseminated|metastatic cancer_C1384494
C1384494|T047|ca mediastatic|metastatic cancer_C1384494
C1384494|T047|ca met|metastatic cancer_C1384494
C1384494|T047|ca metastases|metastatic cancer_C1384494
C1384494|T047|ca metastasis|metastatic cancer_C1384494
C1384494|T047|metastasis ca|metastatic cancer_C1384494
C1384494|T047|metastatic malignancy|metastatic cancer_C1384494
C1384494|T047|metastasis cancer|metastatic cancer_C1384494
C1384494|T047|metastasis carc|metastatic cancer_C1384494
C1384494|T047|ca metastatic|metastatic cancer_C1384494
C1384494|T047|metastasis carcinoma|metastatic cancer_C1384494
C1384494|T047|metastasis malig|metastatic cancer_C1384494
C1384494|T047|metastasis malignancy|metastatic cancer_C1384494
C1384494|T047|metastasis tumor|metastatic cancer_C1384494
C1384494|T047|ca metastasize|metastatic cancer_C1384494
C1384494|T047|metastases ca|metastatic cancer_C1384494
C1384494|T047|spread adenoca|metastatic cancer_C1384494
C1384494|T047|spread adenocarc|metastatic cancer_C1384494
C1384494|T047|adenocarc metastatic|metastatic cancer_C1384494
C1384494|T047|metastatic carcinoma|metastatic cancer_C1384494
C1384494|T047|spread malig|metastatic cancer_C1384494
C1384494|T047|disseminated adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|spread malignancy|metastatic cancer_C1384494
C1384494|T047|disseminated adenocarc|metastatic cancer_C1384494
C1384494|T047|spread tumor|metastatic cancer_C1384494
C1384494|T047|disseminated adenoca|metastatic cancer_C1384494
C1384494|T047|carc spread|metastatic cancer_C1384494
C1384494|T047|tumor disseminated|metastatic cancer_C1384494
C1384494|T047|carcinoma disseminated|metastatic cancer_C1384494
C1384494|T047|mediastatic tumor|metastatic cancer_C1384494
C1384494|T047|carcinoma mediastatic|metastatic cancer_C1384494
C1384494|T047|carcinoma met|metastatic cancer_C1384494
C1384494|T047|adenocarc metastasize|metastatic cancer_C1384494
C1384494|T047|carcinoma metastases|metastatic cancer_C1384494
C1384494|T047|carcinoma metastasize|metastatic cancer_C1384494
C1384494|T047|carcinoma metastatic|metastatic cancer_C1384494
C1384494|T047|tumor mediastatic|metastatic cancer_C1384494
C1384494|T047|tumor met|metastatic cancer_C1384494
C1384494|T047|tumor metastases|metastatic cancer_C1384494
C1384494|T047|tumor metastasis|metastatic cancer_C1384494
C1384494|T047|tumor metastasize|metastatic cancer_C1384494
C1384494|T047|tumor metastatic|metastatic cancer_C1384494
C1384494|T047|mediastatic malignancy|metastatic cancer_C1384494
C1384494|T047|mediastatic malig|metastatic cancer_C1384494
C1384494|T047|malig spread|metastatic cancer_C1384494
C1384494|T047|malignancy disseminated|metastatic cancer_C1384494
C1384494|T047|malignancy mediastatic|metastatic cancer_C1384494
C1384494|T047|mediastatic carcinoma|metastatic cancer_C1384494
C1384494|T047|carcinoma metastasis|metastatic cancer_C1384494
C1384494|T047|adenocarc metastasis|metastatic cancer_C1384494
C1384494|T047|adenocarc metastases|metastatic cancer_C1384494
C1384494|T047|metastatic cancer|metastatic cancer_C1384494
C1384494|T047|metastatic adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|metastatic adenocarc|metastatic cancer_C1384494
C1384494|T047|metastases adenocarc|metastatic cancer_C1384494
C1384494|T047|metastatic adenoca|metastatic cancer_C1384494
C1384494|T047|met carcinoma|metastatic cancer_C1384494
C1384494|T047|met carc|metastatic cancer_C1384494
C1384494|T047|metastatic ca|metastatic cancer_C1384494
C1384494|T047|met cancer|metastatic cancer_C1384494
C1384494|T047|metastatic tumor|metastatic cancer_C1384494
C1384494|T047|met ca|metastatic cancer_C1384494
C1384494|T047|met adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|met adenocarc|metastatic cancer_C1384494
C1384494|T047|met adenoca|metastatic cancer_C1384494
C1384494|T047|spread adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|metastases adenocarcinoma|metastatic cancer_C1384494
C1384494|T047|adenocarc met|metastatic cancer_C1384494
C1384494|T047|adenoca mediastatic|metastatic cancer_C1384494
C1384494|T047|metastases adenoca|metastatic cancer_C1384494
C1384494|T047|adenocarc mediastatic|metastatic cancer_C1384494
C1384494|T047|adenocarc disseminated|metastatic cancer_C1384494
C1384494|T047|adenoca spread|metastatic cancer_C1384494
C1384494|T047|disseminated ca|metastatic cancer_C1384494
C1384494|T047|met malig|metastatic cancer_C1384494
C1384494|T047|disseminated cancer|metastatic cancer_C1384494
C1384494|T047|metastatic carc|metastatic cancer_C1384494
C1384494|T047|met malignancy|metastatic cancer_C1384494
C1384494|T047|disseminated carc|metastatic cancer_C1384494
C1384494|T047|spread carc|metastatic cancer_C1384494
C1384494|T047|spread cancer|metastatic cancer_C1384494
C1384494|T047|met tumor|metastatic cancer_C1384494
C1384494|T047|disseminated carcinoma|metastatic cancer_C1384494
C1384494|T047|spread ca|metastatic cancer_C1384494
C1384494|T047|spread carcinoma|metastatic cancer_C1384494
C2348819|T033|Triple Negative|Triple Negative_C2348819
